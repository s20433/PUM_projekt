��~      �!sklearn.neighbors._classification��KNeighborsClassifier���)��}�(�n_neighbors�K�radius�N�	algorithm��auto��	leaf_size�K�metric��	minkowski��metric_params�N�p�K�n_jobs�N�weights��uniform��n_features_in_�K9�outputs_2d_���classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C                              �t�b�_y�hhK ��h��R�(KM@��h �i4�����R�(Kh$NNNJ����J����K t�b�B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �t�b�effective_metric_params_�}��effective_metric_��	euclidean��_fit_method��brute��_fit_X�hhK ��h��R�(KM@K9��h �f4�����R�(Kh$NNNJ����J����K t�b�B  �Λ�k�;���#?�q��[;]n�?n_m����>�	���C?��|2@G�@�༳�Ŀ����e�U�4�LF?j���%P���ᶾ���>��'���S?�R��q�>,��T	w>gQn��ن?�겿�B�?F�̿;�?R�ۿ<�*=䏿lJ�8�c����!?����lS7?D��H�>���C�>��?�z�?���=?>?{g�?M�����y"��k�?�U�
�����?���?kMY?��?��>-��>�z���mn?c��>�n�>��žiK!@��<?R`6��S:>�E�_��N��?��e����>�m>��	�(�ֿv���'�=T�&��JE�gQ�އ�?�3>KZ?�x�?��u@�'@-��@Oh�@�f�@�L�@���@»�@�{�>h�@�F��3@�Q��/>ژ�>E�,@�Y�=�?�@`�L?�쎿{:?ꢄ�ɯ?�6���ϼ�Ⱦlg��t��+�9����?�g��{�?�w8�(�6�P�A?(뷾R��:�ľ�D��z?z9X?3 ?>�v<?�5Ծ�R�@Ǟ
?!�&@�<��4@
��?���?���?!��?���?De�u�:?R��>~�>�*�=�2�1)��K�>��Ⱦ�� ��7�C�l>AW�?�\��)/��:w��@E���ӿ��(�z�!?�������,>��?XJ5>e
Ͼ�G�;6��`=���=���О����۝��/�>�"�>�W$�i��S]�>��b� �
?!�(��0>�<���ρ���/?�?5Y<>�h޿l�H�GN�>z���<���>�3�>u�.����������i��k9��A�<Ҵr�I�����i��U����S�#7�?�$k=;����Ջ>��@l��>�9>�g>�A(@�_Y��ᕾ�-?��v?��)���,����>tl��q?��)�P��=�d]�lb�>�T�=�?(��?w	?�xf>6���t?٤�?�>R��R���"�����)1�'����^D�����t�ɽ��q��՗��<�>�>w1����̾.�?��4�Е�?\����Z&@
����?G�,@*���]�?η����?n�/��>��S�y�6?!��>��>���J�?����Io�]=����6?d�s�����Ԥ>S�=2Zl>���=��P>j;�=4�K?lGO?,̎�Ц���Q���:���=>�س>�4�zj�[`>Z�w�2�R��S?�zJ�JJ�?��2���>��X�H�m>���?6z=�X����V<��k��Ȭ����Uɿ�|�>���ۨ?Vl��#d1?X������">hӽ&�7>��&?�@I?�?}�> ��?	I?��A?��v?�f�>�V&���$?q�u���F��	�[�>i@���=��>��/�H]���=U�>�y$�Sy?k�:?�w?�1؜�k4)��W?y��;e�=� D�[�w>�\?��\����=kd����>?GѪ=���|�%?An}��pt��	������gžWT=qw��?0�Ѿ
me>9ιN���ߘ>�(�>-$�>���=f�1�
?�ʹ��x� 77���=P⾴� �X3¿ʅ�?��2@!�@�y?(�H?0�?hf>�բ?��6>[����������>c�@|P��M���y����=o���ޕw?E��?SRǾ���=�[נ�N<�B뫿��L�^��?PQ#@;��?��@L��@�2@;Á@Te�@|�e@e��@K�K>��@�I�<2pY?��>̀/�Y?D�C@4΋?��a@�V�?N��?�?�@éH�����T�C��/@���v����־��������܉!=?�<��;+?������>��>��;>�-T>Cg��+5�����&��RO?w�ᥦ>2BI�.��>��{�"+1�M`�Q��?�b3�f�3�K�k����>��h��Cr��m�,��������?�H�S(W��=���,�;E�ˑ���~��B�=�g?��H����$�d?����b�(�����yi?�ь�Q��v�x�EՁ?�Ⓙꢄ��Ο?�]��	N�?	؛>��x��-�������u��Ǘ�^}���e���e�C�ؾL]�?e�>>��q=08)>&�-�
��>�JU�L���H�پ#��? �I>CS>�����>ڝ\>�Z?�E��%�E�Ͼ�c�� t<J�ſw�m��B���ъ�~�Q�lZ��/N�H�����j?��>Z�>wx=���>׺Ѿ�
2��2�e?ޠ��ٷ;?�H?F��?�CC?ꢄ��'�꘩���ܽI���Fo��3rB=$9�`�;�ãƿۥӾB��� ��O:�>�Ჾ�����a�>Y��
o�kc�?�
?0�B`�>�R;?9�>����#k�?]7h>
�>���u�F?�Ͷ>�!���Q�ߥ��.�?�(@��n?(�>�,G??��?��?!�B�M�Q�@Ğ>lFV>U��=騿����UE�Еn�����VT��0	?���m��;�ؾ�U���%����?`3���D3�T@�?��8��}@}V�M^C@�$���a��ݓ���;Q�De׼i2�>����iz?_�?9k@U{�>��2?������>u�><�[��	�<D5��@�E�՟2��j�������=YK4����	� ���F>��<���ο��=%B�h�>���|䉾JKž��>�C�>�ґ>4�\?�C�?�%z?��?6$G>!I�?� ��;�?�U�a1�%E=����8D?e�>?o{��em?��W��X9?������n?T�p?&�
?��뾬h�� �:g?`��ݚ�
vڽ��>��J�X���>4�>��>������]�3C�����>nd3�<ݩ��|!��	��摾3o���A��+2P����>5��"��:��.���)����;V"���>���>�Ծ�~��`O�N� ?�>>����
?�>K?$�?���UT����>sL/�#�>:泿fj@�.�~�[N�>E�����˼����y���5>'Y���>
s��1i�Sz ?Т�?�EH����|��>������"�>�=����,�޾���pO�|!?��"��e}?X���>�u�@��҅��*�ھ8w��W�?Q�>n���
Ui�l�V>˼z-��f?�!���?#�0�`�@!�6��X�֨�?~򘾄�>`x>\��"�K�ǂ2�Ҙ?<�;>դI?�/K?��?}D9?V�?�i?6]�>f*��V>�`a��<��]M�!uz=_�𾻮o?c~�S���g�?h-��(�e>��;>�q?�;���]X^��XQ=��м�Pο�C���l�?��Ž�!��ZR�Xy�?�3�=�P>'J���.�?V��\R�>�I��S�g�^��>o.����<��f�=��>����3�>U���R����������S��>�q<q u���h?��5?�T�>v}?z� ?�]@?Z�?ޙ�?��>����&HV?-)?!c=����Hu?��>��1?:��>�It?j)=>ݾ,>�z߾��>�;�?�ߟ��̷�J�4>J?5\��[�8��n�����\�>��ſW�>=f�_�d�?�h�R�W>��7��J?���l6i?L쳿���?دM�9�>�m�.��A��M�0?��H?�@@��[�?C�2?}S����ž|L���r�U�����g���M���胰?Ƒ�?�;��+W;b>vF���4>�p	=��<F�?D(�?-ݽG���˯?�\�"�b?j�8�JZ~>������<|��Y��I��N^�?�Z�q1F=N0���:�='�%��ڣ��
%��Y�?�4��VsV>�YL�*A�>5o(�:蕾\坿��?_Ő=_N@�Җ��
?P��k?q�>�b�؉�?jݾ7��?�0��>�?����"32?�G6?x��=��"�v�о�b>�Ĕ?�F���t��e��I�?�C�0���Щ��h ?�׾p��V�پ;���|�S����A�¾i���:���}̾qH���,����=d��閾F�����j>�J�=Jv��R���-<\��>.ڐ�nf��M���C?�-*�B�A�{�X��r?��Ǿ�B\@��>�4?������?�0�.�	?#(!�l�>ba(�:�?��࿘K迿v���>��!?�����^����?��@"l�>Z�?�Z�?��?����5@��V?z��?�iM���@��>s��?�t�>���?���9ʯ?A�j>k��?#���3�?oŶ?��c?�����?(½?�>"j��h��>H�@��>ɬ~��W�>ް@C�@K|�+^�?b��%2��8@�<�?Q\@RÛ�юH?<�����m��y��>z"o�y�o�ˊտ�P�?�q0����?o����=��1?�}?��'��4���\ =�����-��5�}�-*�%�==y�G��?��s�ܑ?No�>D/�@�z�?5�@|��?�k@���?�*?f~?��m?@��;���=rp3�w@�=#�.&"?K#s=�!@�=�\&@�G:�<6a�R&��6[�>�
?{�?�I3�k�ʼE�D�hzM�%�&�� o��־��j���������m���짩�J�G?	�>�;?���`?�A$�c��dzO���m���:%o��6���q����y瀿�&�=�Z���?�j�>1@>3� �
`??�1!��2�;�.��- ?��.�����9�}�\��OӾI�?������6I�G?��������@�������?"��>|����&��Fv�ٞ��`��+�>
�>��xu�G'>"T?�x�?/�?=t#>�pz��QK�5��2�Ⱦ2W?3� ���<��[���f�fE�3>�<��ľ���?1�T?�ʫ>W�{?}W ?ߊ�� ��>X[���T?��	[�5ѹ����>�zȿJ`�>*�6��(�5*=����=>OD�)��?�,?1ھ�����?�l?NQ��������R?`��=�䱿L����y�>f�<���e���_?�������>[�O�.�?��m�״�?`=�?����1�`�2�ш=f{?�F����N�G���>��H�?<��ۉP?M� ?��>\ʾ��>�:Ͼ�2@?r3���!��U#�K��>KΊ��T�>z�*����?:��<���>K�ݾ|�?~b�;K���J�`qo�Ǽ8�B�S��ܽ&?�I�-Fƾ7�2�?J1-�sS�>����Z��$B��)��Y/?��{>�!5?�*?�2?QĢ>,k�>xp�> =\�Y�W��Љe>ͦ�>�B?>_���|I>�<G?�&�=����0�"���6��p0��LѾ*�-�辑=���B�Iѐ�\J �?�a�A<t��ה>a8-�j�0>����y�>O\��Z?LQD��j->s3�k@�?W͠��0���>�}�n?sTN���Á���>�5�ꢄ�,/>�D?ƙ?��'>�f�>w��6�0?��#?��6�>�����n�'��?�d?~�e?��?�� ��*z�h"־/B<>���������>�⡾�k��d���@?V��D�F@�w?��>�ˮ?-f����?x�0?\�{_+?gX�Ms'>���q�>�%^?i5>��뿝�2?S����@�l�>3t!?&R@�*�>~y�0���d�?��4?�
?���?m�����?��W?m�1��QV?�O���?g3�@��?	���#����	���?�h�?Wgh=���z�>b#+��#>�$w�T�Y>��>5��?N�@��@x��u�Q?5�-@L0�><%�>䨑?%i�?A���cp?}'�=�c"�K�<�y�� VZ��dS�סE��,,�(@����a�E�	�=I:}�q�+��8q>N�{�K��އ:�� �>/4����v??c?��6��+�?1Ž9��������-?ˡv�W�G�6HX�{r������&�<�: �>fE�?���?%�v?����~>����iq?\L޽��>K�k�o��?�ZB>Pp���:	�"�?�7�X�����W�a�?g-m���>��`+���y��r�c$G���J�.G>��s�!?�G���>y���
~>�~v�w鐾�A���v?���a���ᾄM��$ >(?��U�n����ؾ�8�S6��Y��?&�����?�]���i�?^<�q9�?W~�?aJ���D�,���k�-?F�K�(Ď���W��C�?Zԉ>��I��6�L�?�H����{����b��~�˾O8���1�E��$�#�>*+>����]=1��'�N�繿ɏ��Y>�8	�f̏�2����>��ؾ�\ƿye���q?�����E��	�>��?���?�)��愊�� �?�%Z?�@#@6�W?���?.��>>?��c?t\�?9�.>�G>��)��A�?���ټ�>С�=�@�$h����?�K�=10>P�.����?G&���a>V�&?��0?͢�;�?���?��?��B>���>&,?9������[J?a�2��X��g��L�=�z='à�F?�:*U?>~�?���?��?<&/>�aw����?�� �.ꑿ,���
?���t�>�Կ����׀=��+�u�,�I_�;zb,���?�x�?��>������e���O�4@u�B�"��>Ѕ�]��Y���I��J{ľtj��>���?;��۷��t�)�↿�ʾ�:��4P�����1>�( �� �>Z��Ĭ|�,Կ�m$���#���>`�տ�Y@���>�ѳ>�=���>�L8?QXv?�b��׀?�=>�� @ꢄ����?�	�����=�Yu��dC?^��� a?,ن�n>?N����aվ1�̾n8���\���	>�.��S�?�p�y�ܾf7���?�>y�q�qm���%4�8�Z>���hʉ�����*4�<�ܽ�d"��g}���>�����G ?vr�k >x1���?[V��h�>����c'�?@W�~Ĥ>�^ÿ�Т?�揿۵�.��)�?k��Wؾg�ƿ�B?<���sS�>xݺ����?����i��G0�384?$  �f�q>�`[�P��??����ɛ���>����������7)��}`?���>փ�>�T*>`��T]A=��?��A>/�:�9콞�����?�n��z�E?����K(?M�O?�~�?�>��y?z��>��7��N�Y�>�ɦ? XZ=!��>��0?(X�4�?h� ?P�l?#M%@�� ?��?n��>��?w��>��?��H?\=�?���	v>�]D�e��
���.*����+ٶ�k ��KȾ�达{�=Y�"�+k$�8D?��>�MI���4?�g�	k*���k�`��?�u
�	ᙿ�c ���@W������#���/E?�����l�(�2{m>��D�����\�i�>�0��	�>�R���e<A�0��m??)�������()�>���Gff�<�>�5b?�����]��|�1��U�8$ÿ�	.?o_���>������c��11��^��O���3�Q/���擿|���5����>R	�m�پٕ�v��?kaf�d͎�B�5��s��)f���þ4}T�9�Ͽ��f��棾���'Ξ�\m�����0~,���w�q0p�[���r���7M���@���M>��<�(�?�x����8?d6`�r��?����[���,����^�%ľ(
�m��|J��
��U��
>K���L�]?�6۾
��>�eB�*��>!��W�>�쾉(�=�~>������<��?7�?�k�?ȟ��h׾RW���?-;�>�\*?��&�~U!?-T^>������a��	��Z+�?�-̾�%=7���!?%s]���%��O��F�=MK�N��>��:��꿾mD��l�� ��a�S����>iQ?P��59�+8?�C�R<���`�a�?�P��U���7�M�?�=?��9@9�>�����sC�i؅?v��ye�=Q��<�UQ=��>��?���>9ܾ��g��;�?��>U�J�v�����?��2?��e>�Z�$�#��庾�@�*ƿ�J�?�X�\s@��r	@�����	@����R�=�	_>���?.>�߷>�]+>�E�?��%?�]��Ǒ����>�(�;z�?�)ʿ��?�P�?\p@/�=��@��v?�h����?SÖ��	��JL2?ܼ?}}?2�Ͼ�?����;a�?P��?��־ir~�h��>:�
�In2?}]��b�=�G�>־�>��z����?�%e�x�>�ѿ��@*���jȻ?����C8�?�}�� ��?�A?�*VY?g�'>�#?�c0?m�?�>��?�S�>�f2?������?0P����?�i��\{?�,<��4?u�T�l��>�>L>ܖ��|�������G=	ľ�
d�U2�>�����?w�.�ߡ�>��羫{f?�h?P�><�6�2��=c(�>rj=?�l�X�ȽƜy���>?��<��nɾ��W�;z-�g���!�3V����<#��AɆ�$�Ӿ���<b�=+����qs>�Y��iX��O#���Ⱦn�^�9�i�����(U���<��a>/��9��Nt�>Yf��e�ؾ�]��ov�>\�0���>� =>���	D���\s��`��i^����� �l��J��π�R�<41=�`�=�t���*���*���)h�<�w��(@������
����+�/@�x�g\d�������?te4�5r��r[��x�?�)��z҂��c���4� K�ya�?�24�|QֿP����?B@N��@l��.�=~�@eqU?�=r�-"��_i@��쾛�D�RJ>�k�8@�f>�ȿ�����Λ�Z�Y���6�e׺�V�i>�y'?2u�?�2<?�&�?�#3?��@(؎?[�?>�>�_�F���=?��O?�s%@�ۼ�	.?��7?R�O�����0�t�9%�>r*��U�Y����N��>qÓ�ʫm�F_C����)����\�iF�g�Δ<���=�C���7?��@�.�?���I��>M�;����"���3>�
'��$?�p1���=�'Ž�)>�ʑN��U��~?P}��p焿v�>"�������?0x��䝾��B�i�ľ^������uw��I=>�s�q��������>[�2�#%�>Ϡξ=|�?<����r�=�^>�(?��8�^4c���5?��>���Ɍg�|�s?*$�>�̂�U;����>\_�����$M�[`C�5��@����>��d׈>Q��al9?-%;��[�>싾̂�?�F�>>4�B?w6�;�z���H?H��?��
�Z���7 �)x>�p���X�T�h���^�����>�B�?5�=M �?b��?�[�>J��>@�������֕�ֿ���@�=�5��c뢿]�]�V=�*���ܽ�,YV�`?��V���.Ľ�A��Q|?�a¾�Θ?��>�5@�l^<=�@+�F>N	�?�?VԿ>����B~�	]׽�)���4�½��_r�>"L���U�o��<@��?�M}?K�þ�2�?cM�qɠ?��l��/?Xr��\���?� �?Ű�.xz��m>��c�>Y�>�X�?�͍�j�:?C�?�^���)�~}�?N�	?�t�>�п�r?@�Ԫ?���?����?��@`��?�K�?��@�B@�@r�4@��`@���?�"�?�G�?��?Z����G>!߂?l��>K���U�3�/�@ܛ?�>ӿau�=|��g_���#���ٽ,����±?B��=�҅?M��y�?�r^��n�?~�?����X־��?�I�>L+�?�*�����}tɾ�q�=o7�>B���7P�>0�=��Y>�8�����>��%��ǉ?H�d��>$�M�MI1�mT¾�?��)	{����<�&����#?�EO�{{��v�Ҿ�+�?�,�w�ξo�>�����Oa��"�SP+>w���}x6���m?wx�>�
?�(2��}������Ň��r�?=zF�s�?���9�?�	>����?���?޲<�ο�����¿
s���c��'n�ls�� ^>?��V�"�>�!�H9=�����Ǳ>ϴ��,��������?KB��W#ÿ��g�� �>	4�� ������?,��;�QX��U��Q?��`�{=��]�ƍ�>���ױ���B����l��?�`���#����=}����U���#����?�nྩd�?���$�?������</�`��?c�"?E'?͹D��M�>�G;�]-�@�<�>���ӓ?��̿�T�?`:�?)
/@;�ξ���@�,s?�nh?�Q�����?��>�4J@����Z�@��)?�@y�>l$�?�W4?3I@"+�?7?R@wپp�C@���?cN>@z6
��ٴ@Я�?=�I@���-<n?�)?��-@/_��<�?�U��>�'�� ������,�>�hž7]?b��Q!?��W�Th½����=j�{��	~E��o��V���V�fG=& ���?�`c�6�Ҿp\���:@>]b8��i��ǣ�e������4��j���	eھ���n>��宾c"�>��Z�a�?�8�Pr>?�-l�R��?��7�:ϑ>�#�4\?g�8�_!��c#��t~?kmi��t/�7���4�>8�_��U�*2F?�j?�1ҿ�Ͼ^%m�~��?RJt����;��;	�3?ny��"d� G9?��e���Duʿ��F����?˳,��U@��)����?6�n>��F@
�����?WE`?�]�?�����?كh?���>��۾���>	ћ?1�]���{���o>v�w?.�=M��>��g?a]?���?}��?Z"�? ��?[@0��?��?:X�>�C�?�Q�?pG�?� �>Wj�?�U��H>?c��D�H�\����"�?��	\�?�&ܾ��?ag�>D��>�[��\ɿ�X�>:��Y�1����>��*?���?~�ɾ6��?a=ݾ�<V?UW>p��=�~T��Y%> {N��;Q��l�>e����žQ}!���3^����w
)��g��ޤǾ��XW���V�c��Gŝ��M�|CA�4U��r�=_x���%�~��a><��=�U��;���x?��
@�U=w���25ڼ	Q�<렾�ƾd���v̹�}&��a�>M�@��E���?:h�?	���	A�~��>��8�7�*�<���;�Q>���?�r#���?�,����f@r�7?�@�>?���?3_��j!�aK��k��k���S�^�R4�?�K�>�-ڽ���<��޿��#��d�����{(?�_`=�k�?��6��(���Z���?�����H?�M�?����j�?Ld!��l�=��-�ڸ>l�f��Ƚ��a����t/��%-?��?�I�>�|��W7?�BG�̐���}N��A\�:�L� )+?�>��At?e�($¾?�Y�O?C^}�ى��Nd��|L?��.�_� ?� 4�V]x?9�@�e�?�F��$�?$�n��;�?�9a���[?"���St?�4D�C��)�W��?"d�����*'���?����w6�;�Dz�2��?�@��S@`�>O��?aqO?ҭ@�?���?�H��B�P����/@3���� @)m ?�?>�B�(�?`^(>$dV?ٯ��،?a��?���?h;�=d>[�$@���?���?g$�?�/C@<3@m?��K?O�.�6�`>v^����:?����� d��\?��/?���>F�?L"���J��3q������)ɾ�
���ߘ����������v?	XD?+��%R��?E&����?�~:����?K�C���?��|�k��>b��>�$��s���Z��v2����=9%z�	o̿a~�@`�?����fɼ�/���p�?#`�q��>��l�-
~>+J��)�>�9g�OFW?o����k>�hz��ƒ?J)��3�?��:���?�ڕ��9�>��[��q���'Z��ށ?r�O��:Ƚ/�&���9?d#&��f��U?v5Y?�u��� �<;K?�|=�^����>��ʾB�?�������|���)��F���e煿��}���V�?�>�.*��D���P�-մ>x7�?�ݓ��"��{��?�P~>�p���B>���?��=����L�?�B?>H]��rU>ȁ�?wt@?,�M?�(+����?P��>�
@6	>��?$l?O�
@ygF>�% �^�G���?t�h>�\��6$Z?���?>�$?)_M�����sS�>S�$?	U�h�t�}��>K8?fvE����>�J���?>,#�� �>%�>V� �Zo�)8<=�-�^ ѽ3��C��f����;'|�s�'�C_>�����쾤�����?JiX>���>�P�N�$�>�c^>o�Z>d��=�QR���\=�|�մ���K��������T�fY������>~�/�ۀ	��0�1�a?�w�=MV߽� ���>�:E��U���ѽV���> q���ށ>:��{��?;!C���?TX�c���������콲�!�V�j=�pp?]~�?#c��.u?3��g�@�q�N���Y�����?]����G���6���K}?�Y������K�n�%??�6�a���~��v����"U��Z�.v��s����h�g�#g�/�j�[�����?��a�c���2S�t?dx�ɂ��ч�c�>��Q��}�?���?�iٿo��>r��Z���<{������P��$Ai��:���p�����<�7>�痾��s?G��?} Q?�r��ro�?l;����*�V�n�?T��e;����c�&=�?�/"�X���]f���޾����hU��YZ[�%���؃�	�>�,�����w��*�2?�H��gXڿ}�y�Ɣ�>����&w�����G��?$���)+'�2~�]#�?J	���{1��֑��U�8��Ŷ�?���|V?�1[���V?t�=J�=?�B2�H?@�X&���#��W��>a���>��t�0���u�?�&�?��8��?e~==.�ߧK@���<Y�;��Rʿ/��?�K5>^$$>�h%��ڡ=����_�z<����v��?tZP�t`ͽ��P�Mt�<G_���>�yܾ�>���܏�=������ ?w�-�n�|?(վ�?�5����>��>�{?sS�>ڙ�?qz��h�?��?K��?e�;?T�?&��>1��?&�?\d�>� ?f�>e�?�T6�K@&��?�!>��U?��>�@������%��7@ozξ����fU���>OvO�i5�>Jy�ԅ�?�_��� ?��ɾ�� ?�j��Gs����X>����>��A>��>�m�"���)�vx,�l�������wI��V����/-7�.�"?�10��U�)�L��a�$��?㹝�$��>��G�]��?6��&08?#
��p�ԾL4̾cs�=�ŗ��=*�.@@���-�'��؀�,X�?��7��˾��'��>�4�ʐ��Ý�{��?V`p�A�P�t�.�?���� J�>�n�0	s>C1g�۾��=7U��4���m��_��Y;��,A�sJ�,�˾�;K�,9����=�Ӿ�����x�9���d0þ�␿�� �Ev<�P�0�z�-�|\>bp����'�L(�����z@��%��YW=�dv=���=f���>��>�$6ž���b�X?���V��HfX�1-B?򬾶�z?���=�q�;�D��ʚ�X�j��?�A���`�?�` ?��5�;�URB��>H��> ���-�?eH&?��޿N�0�VH����>�=�>�0׾�eT�Wn?`xa��C���>��L�A�<I龄�>~;�>�zf�q>�У���d�ꤾ�� N��m*�.�;����C@_�U�ξ���b>�γ>�ހ=^���xS?-Y���� ��c�H��?Ԙi�w(���ܾ���?i۽�������>N��<K`뾲Nп��}>	 ��~����5�����?���x/���?�U��Zн�.P���?s�U�jP�ep�S�@�����!��V�����?�$������eQ=�� ��O���c�����J��O?����y�3�_8�
o�>+���c�?C��?���`��3X�����k��=�{ѽuY��V�S+�Dej�Š]�؉��� �?�4�?[�p�H�п�D?=�<?6�P�4��k3*?��j>d��ͼN=����k\���־�̓��$�=�fѾ]�>�3�=j�k>�ܾ�E�>pr��p�6�?�Ҿ��]>�ھ�j_<�
 �v�?b��t����?�%-���?����/z?V�࿹�׽�?����>28���G�[�>� ��ó�V�|��鿌g&��?Х�?rK��@��>��?�?�W��M[�?�C?ϑ�@�+m�Oa�?CA��.@HC޿q�?k0��t��?�y'���?����c�?i+%?��?����|�?���?U�a?�����>ql�?�l�?�|����Z@�J�??@O䗿��@�� �,T��/�?�~!�ͪ�?����o=#�&��/9?�-���.?���������>�5;c
������.A�{&@0�@9��?���e.�@���>�
I? ��>�l�?�6$��m@ݬ4�M
�?�o��!T@K�&>O�?o���$#@���U.@�6��ו�?�>�s7,?�M��,�>Ä ?r�_?ke>��V@I��?�@��d���]@��?���?w����?�U���Q?@�Q�π��N�=��T��w���K�>h���K,Z>-�H��OG�	|I>��߾�������>��&�d�-?2�?r���x)���n?��?�$�>e�R>��?���>�َ>��A���|>��>N$?mG0���#�I��:>TWo>��+?s>˿FI�>��%����Kܔ��U��[�K��=
�4����=�����곿}���7�:^�=A爿a�w�����\��?G��?�(@5Pξ�P?-�>w�%?0�E���?&���இ�pV*�Y��?�q�?�v^�4���t?>x��^@�G�>��Ҽ�p���NQ@a��> ��<�� ��!��U��n������G��h��(Y�=1[���W��e��?�8&�ϯ�?��(@r�'@\��@�8@�dA��!@�D�@���?��#@����5#?������?
����%?]M�?hخ?4`���l�>N��?T�)��%?�����	2?������>�P���gI��Y3��N�>�;�>*���?3>t,)?Piƾ��M����.}w?�m�~�*? �p��!�>_!��!�=[[�CɃ?{m�����
�~ņ?�U�����>�9ž��?i���hH)?�0�����>��=�O�>a{�����>�#����?f��>��A��'����>����	��]x:=�?B>?4`����?=��MP�z�� н�����&�>(-ǽ���oE��z�[�Q|[�?~$��<�[b��Z#���j���	��b�>�T��3~?\��򲫽������I?�����C�i1G��l�>�S��Q7%�υ��+��~ɼ���C�=Ը>�WV?W�-�l�ɽ`�5���>�C2�4P���~c�J��A�"?m�&>�r�>����l�u?ȫ��H���:s�-�?X�M>�U���?�D��,�N�<y����?⭔��K�?�]���?9u��Ě?�9�?�25>����.��1T��1Jl?.�s�`���wf���O-?�k��~0�qc[�R#�?lB���ݾ����E?j� ��T�>�3v���>������<���������T�X�>�=U��7�r^J��
U?�P��E�;� ��q?6F�����R����?��1��tt���!�z?��(�ꢄ��H>j(??y�?)��>�/�=z¾֪�?[���z:?�޷�S迿~�Ŀ����N�?|�?������=C�����u�_�����?OH;>b���
��O�?ޕ�ѱ"�UA��gD?�'S�z�:�U��ȧ��۾ZP����׾?g��6���\(��J>M��FS#?�%@dT@�Ő?dmB@��@��@�8�>�?G�?2�(vr��n��
�?��d�h;ľ� >�:�?��%�Cۀ?4����?4E���O�>떿��s?����#�[}�>�{�>|r��e[j��2 ����?��?���3?mZ4�7V�?��?fJ�?66�?釦?y�?S@O4��Ӹ�?�yx?�=�?P��C�S?��N?G�@�ZC�q�?4(���#?/R2��L�?h
�㿫?�&�>��9@o�8��,\@���?��@�����@�?��@E����T@�� �]hȾ���?[?��l?�h>u{�>���>�zԽ���>�}�ڏ>��Y(��žR�t?��R?{Ŋ���*��6׾���r!>w��>ٌ�)�Ž#�>j��>v�>���>��>�x.?>� i?��h>�@� �?Y��?v|�?��@ؼA@��h����>�c��.i*>>/���&?�v����?@�>sX���p�?�?#�?�@>�+=��;��?.>��3��
?���v��?�˽���?�:@�Kʾ ??p'+�B��?)�h���Q@ CD@P����>�,A>0�羑��>
|?����I<���<�'?�W�=�,��솧�O�>:�(�t��?�翰uo>�"?��s?�SA�_�0?�Z�?5�?�Z?A^�?���??�!@2%�>��$@�@]>�\@^�H>L�@T�j�]�:?���>������Y�?{�?�&�>������]?�U�����`Ӡ?���:��?>@�@5��?�󘽌��?Ru?r�;?��??);8=D����黁糿�j�ԫ->�V!�V��?�_�?5�0?B[Ƚ�M�>� ?�5>^󂾺?�>X.�>2$�>�P��֚H?�U?b'�?��?��_�N֖?�Pl?,��?�i@?�Hj?�È?z�?�@�?��=?d��?
b�?p�P@lX?��}@5"�?IWf@r ��"@0(�>%'D?�� ��`�Gb?o�=�\@��?5��?��?����-��?�6�>IZ�?B.�?i��>�t�?��=R�C���%��?���'G�>���?ٴ�= ���,��ٺ>]��Z���gɽ��[>�9ܾ`��G���t�=94F>G"V?��t?sIr>���*�>�[�>w���:s�>]��;(@?������5=>�9>�]�����<��?ů?�����?��?]��?�U�����-�;�>;��=���%�?�"��˅?��M����?�����X�?s=�?�q&�������T=�s���?Qc������e�>	J?�.9��KL�x���N��>������L���$"<�'�=�O�=��C���֫��>n�O��d!���D�=� ����dn����>v��>��@��$�:bJ�.��?�������4��EA?�7s���c������>`5&�ꢄ�:]���?��c?y9Y?ck?��h�熥?o��*'�?˞��� ��[F>4�D?��սݯ�?��^?a���(y�6|���p?(�>�=q�pm����?��>'z���ڃ;�:�>��>�F���у=��3>��? �a�^�>,�ͽP�?%�f�C�?7[E��α?�	���?P6���g�?ݽ�/*�?�:��+��>�|?h��g����[�?юU>�U���E�f�%����� ���_�?�NG�D��?�� �Ǟ�?����?l��?P�=����x�,�e ����y?YЂ�6�[��/��#L[>�&P�V>��ߣc��vL?�Z�gE���Qk�P�>��f��̾|���5�<,���+]2���^����̾�6P�M����❿��ï=ľQ�3���P�mu2?=;C�I����	���d?�?�d��=2�<�f?�+���
?v�6��$�?ds�=_��?~�/�g?$V�s�g+���>���l��%#���>*D[?�;��\�&�v�BK�>�v?5&><ɔ?���N8>I�9��=�[?�r8?�{�=�`>7�=,J�?�]��!��>��j��p�>O����?f�߾5P>s�B�骾ﭨ��<?��ʾ��>�t�0�>%���!= >�"P�Q��>�ow���?��D��!�?��v?��	���V>�<e�}�#�U.?���9�p?1>�<Ni?�>F��? k�?
Le=b�b���9�5��?��E���ľ����׾wVX��~#�Z:�D��V(�	ʿ�V)�\��������{���;��ڀ�4D"����>�U=�q?9����?�E9^?��i>@:�?8�?m܈=�r2?��?P.�?��;��:?�?�X�>[���
��W��>� �>|���x�=���>�I���)�;�I�����>y����`?�xĿ�<4?|W��Fn��x�{>j��V(�>�>W���&c?��?��?J˭�0�=�Y�>���>�KM>��t?g骾��4>l�?BP?�����A��h�>"t? f߾�G����?��?s��)��md?���>�ɾ!d�/~>4ee>q�޾��h��~I��W���ľˋ�:���<��2��Xǽ�|��Λ�Uv�}�u<�YN�=���޿���'>Hu�=��?ek��K? �?=ؒ�=1jc>Z���1���!���rE=O�ݾTY?d�l>Q{I>�[߾����o,�)z�?Ak����Z¾��=p�K�3[ �������?���'E���+�/�B<њ)�c�+>��A�cQ�>Ϣ�$��>�������l���>Sq ��$��7hs�o��?i����;]f��?!L���U��ɾ���>�+��5v?� ?Y�)�u??�qp�k�C?�"�\0��U.�<;w?�f �4�x�j�*�]���$�?�۶�=�I��5?���O���@��/��Ͷ-���?�h>��>�}>}���[�̨̿�>ܾ�/�>�����]?��>���?u؅�I?�>CN=~���lw�P��z�ڼ�e�@�?;l?��1?U�V�~Z$?�t����)��E��[-A?��v?�^�>n#(�iI(>�.����>�+o�iA?�g����>�"H���G���?��2>�M5�L�(���?	�Z�x"�M���ʙ?�㋿�\�>:��l4�?��ٸ�����ƴ?v)J�u���Ff8���^>߉��K����v�=��>W�:�|,?9�\�f�>�~��p�x?
���+!?��(�3J�?���Op���T="�k?{[;�(���ѻ�'?2�	���H?�ƿ���?]����#=p��?KA�>m�Z���M?��>�T>z@�� @$��=f�{���=i��e���%@ޒÿ�K?`�n�0�?u !��Js?�����?�V��oG�?T�k���V?��Ͼ� ?���d��?@!7�a%8@�5���L@b�����?�v��;<@�i�f�@�뿄n@��-�\�>@��2��>�e<��Nr?�6���d?5����d?b���M�?x?B.m?:Q�@��y�5&?��>�@i>/צ?N0|��d}�����(�@�>�\�v%����?��@���;=l��>ÏG@�~���?��?��.@o�?�0�@)x�?Qr@�}��*DL@j�o>r}?6�=aN�?�b?���>�ъ?���?ψ>�͕?*X�>�3�?�i�>$5�>��W?as5?�y���(>�k޽P�F?���)M����>�8�>�U���?unR?�i@��9?/�?��?b��?n��>`'@2=�{�@>�Y>�]-���D@Sj6��m�V 4�W��=,�&��o�>)��?��M?_��?p?0�6?�ۖ?�@}/U?Xt?�]�>6#W@��;@@�?��`@o{@O@-=>*�@<�?ͬF@�'Կ�+�>I�N?n6�?g�> p�@��?n%@Z8�?6�@���?`T@~��?�B?�⚿ӆ�y�?��?��?NO,�\`����X� �0�2��\�>�f���'�4�eT��f�o���ڰ>��A�F�"�+�D?K�;=Pi�N3c���>�^��K/?C��8d�)C���K�=5���4_�[����&�M�??/�R(U?La�?�F�?�A??y4?n֜>�F^?ɤ=>��0?�޴>2�?���DS>��$=��p�=T
��I��I�?F���Ɖ>*�L�q_?�U��j�� '?��`���=;]�=;#@�.V�K��?����R?+�������>�5o>)����o�s���~��>Gd�s`�?�rI�z�<
��qU߾���=�h���I��k�N�����Q@�>�p��9�>�Ѿ~%y?W��ЊZ?\�:>�S�?�G@�|֙?��g?ɓ�?��a>Ed�>�U�>@�>8=Fw��/�>��b>�Eq��s�;���(�?K��>b��;�$��	�8@0���č�JD�!�1��i7���M���qs.�U.,���?��?�(@�@@�v?b���E�?h�¾��ŽlK��G�:SK�ƣ�|@c�0B?؄�<m,?ܠ�>�v?_�!��)���O �'�>��X��˕>��V��r�=�Q�uq�?����.z�>۾r�?m	��Ns������ה?���+}�'��W'K?�F���r�fCH�ꢄ��d�Ʋ�>��o�Ժ�� i��O	��"������ݿ Bd��t=u�=�U�>�a��z�fW����$����ʒ��;@��f��b@H����@_����b@ �f�&��?�"/���p>����3��=�Q?�v>�A��7j�;y�*?8��=�$�?�&��;+�?5=�>	�?�[>��C?ʰ�?�j�?��?.;?p��>j?�(�E?a>D��o>~�Io�̖������^?>pz�'*�d���fB�n��5Gؾf�l>��m��Xn�A~u�	(=��>�{��֜V�
�N��B�>�;S�Kd�=1ԾIuk?mP�� �?��нs,�6� �o��Y;��$�=1��þ�q^ƾ�Y�?-V����F?� ���g?wAǾn��>�/ѽ��z?l�4�\�2�hS�=9=�??;���?�"���?	���x�>�%׽��.>�� �n4�zu�?����}�?%�F�T�B?[�����C>3g��c?aA�� ���,_a�k����?GBѾ����K��?��>��?�mj����?��?i����>X>�i�>���?��)>�N�	�?/G��b��?�����N?�S�<�>�F��\�=�#ſn��>����Y�>�c�
����>�i?(F_�:@DGC?'&�?� ƿF��j�8?��>k��Q�	?�
?sV�=���>
�J<$a�,���,b���ǿ�Y�?R�^�Ž㕿��^Ŀji�>�u'�o]�=	�?
�+��≾<d7@�<���z=��?�~G��4���нm�� ����%?˱�=
-?;1�G���W�?d��y
���6	?[����q�>hb����=I�n؆����������nb��g�F�s��9L��ֳ��P*�0C�r��(Y;�ErK�uS��y�?~��?^jU��F߾A�O����%�Msq��)˽f��n��<+=Y&=���Te�������;�� C�EY�>�g߾SAw����@'H[>���>\� �`B�?��Q���ݾ�M��W
?���p�?�񕾽m�>\�L�&��>R�m���ƾ�,�B��>�U�P��@I�&�G��e��Vp�n��Kx����;�s*�(���m��|?H�L���1>�� ��I]>ʜi?�^?� �>���}	?�+�
ّ����`B1=sZ������"��n?/�>���>�=_K ��S�>/[m?I��B�$�?o�����<���T?�J��3Y��2��C"�>/����S�¾���˾�eI��nZ���w�>��Cx�Y�N��	K?�վ	��>Ι�>�{���3�k0��y>�.���>��V���C?%w&?6/>U�Z?h;ľk	@��ܧ�?��P�����g���蚿�c��`����_��Ҏ�8W��2w/��X�?eۥ�~vS>��S? 2���=?:\{�NŶ�ⵉ�R�0?����jo?'����01@�AG�80@Dl���?.3n��7�><��0��><�x���?�v������V�cq?J��������N�������v��數�����<����7Dh�>���^
������pڿ�����B\@~�>�p��#H>�3�q#�>3��?�a�>�J�>Ծ�>I�?��D?mPH?[����e'�5s2�}B"?0]?��>>A�n�2+k?�ë�d߾��O�S�+�Y�?^%��=�����>�7z?2w�=��>���.�]��[z��]��@��g�>�J>����ž�������^��MI������z���j׾�(X�R"��]���rǟ��Mξo<�X)>�j�
Q@��?t�x��(�?�&�?�@7K�?Ħ@jS/?��'@J��>�Ȩ?�{�?��?�t+?H ����?5��?�j9?ׂ��\~��H@9�%?��0?�p�>Mb�?�5���z��>k�<i��>h�l�b{>�V3�.�?����
��u�>�(�>P �="i�=���=��Y?m����N쾵$�=�v?j�ؾ�������^w?��Ҿt��IҾ��?N���U�i/H���J?D��?�j'@!���Q.>%!~�ۥ��)���u��Ψ?ʁ�?Ÿ�?���?��*@��?n��>�M= ��)#�>���@�?�g�>�W}?��Y��x�)�?������?礧���@T�N@-�
@Bss@۞	@B�?x'��a?վ���?zi���"�>�򪿶�ҽ���?$��>΋	���M?bb���3>!�
�i�;�Y?F	?w1_��k�?sS�>0�<T��j���F���X�>�Gi��(�>R�|�g?HR�����>7��>�>>S��8���Bo��Nw�?�@��룾�A�?~�ɾ��?ޟ�j����ξ:�5?�凾\�#���g��K?
i��&Z�bL�|��>z����8?!�>C!�?G�ѽQ���>�:=v[?����������>쬔>`=R�y(+���?���<a�Oe��?����
? {�3n�6��/�1�-%�?Sz�>� �?��0�ڣ�?�����@�� @a�(��b4���p=X$����S?�z���������߅�?�N�	s��aSd��19?�w��j��=������>��r���r?Jþ��>��r����?C�0�{�>��S־���>i�7E��7�����>� ��+ھ���/�b?��'`t�64�dn\?������|�c�žF�`?[<l�4`����r�J�x?��$��{�<���?�f7<�+�?\��*U�?L�ž�7?��;?t%���M���g>vI�|�5>�̕>,Ӵ������͈>-�7���Q�	�����=A�i��.���,뾼���I�<w�?�/��*��a#?>�5>q�>�)��	1�>��=wt�ߡM���>�[�>͘&�G칽��ּ��?���>�<?���?e��?���?^��>ؔ�?�?{��?|��-y��f�>*<����>9�?��T>��k?i'뾛W?A���I��?*}�?���ʂ��~R?�<5?�?>�D��yV�Q����J�>f��}���ǧ�gߑ�ɧ½��ϿoPξ���{���ſ+�����"�`!��$@��1�̿#=�������䶾ƕ��GL5>-Ӿ#�$���nh�>�R�?�Ԯ=�&q<���>�H/?#���/��
g>�0�>hn#��U����>W�V����>��n��ٖ�Ȳ=�>�>�_���I�=eY���+V��($>�p�;#�m�ΰ��?W�Z�����G�d�>$��K��>o��K��?�ie�e�`? 8Q���c?��m��R�>�
�ċ�>��Y��J����1����>w_;��
�q�����Dyپ�E�>� y>Lh���s��1�	�|����ֱ�����H:�h=:)ƿ$n>��>��?�U�����	&@��?"Z�	����H�͟,>�������!f��<x�
=y�\OA�U%�?۵;@�qR�d��>b�U�n����8_?H�^��Y=?�|#�����|⾦���x սE���Om�>�X�����<��?G<�~��?Hs��R�J@X�#?��]@� X?T�t@M�?�@=r?�#6>����*��:�n-;��%�� M��N�3�?��>���?X�H��
?:��?�V��=Qr?0f�4ܿ��{�Ѡ��4�����w�Eb������T�>�[�>����� ?��y?�wl����?Q�G�V��u>~��>�����>w�> �>����?���] ?�&�=`�>��^���=�l�"��y&�F[��YK�y'6��H���zt�A����o�0��&L��s�?��Z����?���T9'?��0���>T僿/p��V3��U�uմ?U�s�?�������W鄿�5[�P�r��)���Z2��9�D�����S��?±6@�&�=��3?I�q�E�?u��R>��u���?(��{�?�u�m>q���j(?��P���'?N��T��>�ce��e���g��C
?c9��{�W>x��ˢ>���f��>e�7١�*u��TU)���=���0q��Z	�>|���	���pL��u��+����X:v�`}@!{@Q��>�}T?��?2�J?0�_�9�F?�	>�h���h�e��>@��N<,3F?<��?�]��¦ſ��?�=S��?��I���>�:?��>}:m���༅��>Ȧ=H�Q�2�T�R��荾S�-�����9�>�>�0x?�d�>�n�?4Ԏ?6�?��?Q�?��?x��?��?��>�J0@��q>�,@�fe�[�?�?>� ����g�>pU@?��	?��?`I@����;o|?\ ��ٶ�?�2���&?q�*?�#�<��?*tr� gl�}�d>�n��(��o��:,�S�7�qS9�'JԾ��(��?(xҾ�G@> �?4�=@2��P��?���U5@�r?�@>6v?w��?����o퓿�����_#�E�k���^�Z���:�?�Qu�M[?�����?KM�J+�>�����@��w6�;����6�?{��?��y?��8�V���ꎾR�>�+s�ڐn��d*�B�'����t��?���>w�־�6�>e��>�+Q��?*��RC�?�����q��4��P_��9<#@�ڿt=�>��2;#R�f����?�t`?�t�?èB?$6p?�?�@��c>��>?�5$�ݱ?����`?m����k>_8Y?��@�*?�A@V^�?��#@/�*?�@sS�>X=??s>[Ϩ?�G?��>]ڼ?p��>�?�~�>'�?�=k>���>Y�?�� ?�$^��eG@V؝?;�>�_?��p�?�k�>��a�E��>�!>T���k��	�>�#;>ʈ�?��0�?>�
�4ϭ>�j%������R:�٫>gM�=F/��z>,F��R6�Qɼ邼��Iǽ�1��
�����L�Ծiy��Em�Z���*�급�� ����>\y����i>�.b���,��3?�r����,?���A(?��`���o?��q?d�����h�zi>�'��?��x��K������P�D?�E;�TԾ=b���n3�r!3�si����$C�|b[�D?˿�m ���$���E��{�$��>����4��>?ݾ�&?:��>��F?l�v�aKO<��?AL�?9�N�2�>\'9���?�� �f�*+�Bo=>񂄿��v?5��=h�@�"?����^����6?3?6\�m��=��X��vf�וf�rѱ��::=�)@��>w�}?�o�$��>n\��?o��qQ�=���v��?���@�/݇�d�8?)p`�������	y�>I���¾O)���|�>����o��o�Ua�=֨�������y�nT���j��d�>*ҁ��T����o ?�ꖿ�~����c��x�?4���w6�;w�p>B���z�Q��y���lY�P&ֿʔ>����ܧ�@s0>��H>�f��|��5���IW���m���Ծi[�?��^>BKڿ�m?��?Uf���ѿ&x�>!E=���+>4
���>L'?}ԡ<@�>2�̾����2�����Rլ���S�H�f�½�.�~K����=�D?�=��ݿ}�E?@��>�|J>�ܶ���=�<?��V=F�ݿ'-�]�G@#�|?�=l�ƿR{�������?Tt���̳?������?��
��v����=o��Ʋ=�F���y޿5��?:��>��?ʵ?b���4U>Ć�?[>.=�a?�D�>���v?0Ӡ>H��>�l8��ٷ��ž�i�?ZE�p<پV��)b?ۑk�Gs�J{
�s�d>7��`��|�=���;=�?��j@�C2�>�!��{>���G��?7��sS�>sM���+{>�:z?�8�:H�?[љ��Х?�&̾dy�?��M�������ѽ{|ܾ�!=?G"=��>�I�?���R�M����oI?�G�>'����W���4?����l�!������:�>�ѽ4���[�,�r0����𑝾Б<�]�?M%7�k�'?��C�2&��ؾ��Q=�gG����="���,C@�W�:H�?y��N�?�}����A����ͪ�?��7�]�G@���=J� �����������?�<�TOy>84v�|_t>kd��Dn?aap?���=�J�����U7�����<|�`�x�=�_B)�q��pŮ=�1?������sj־U�������諒NH����x��`D��j���<�[p���ؽU�#�`b�����x-���j��ݳ��"��b�Ѿ )p��Đ�����tۿ�`>�a>�(?rj�\��?hD>��?sS�>>�>��/��<�>��8>�+~�f�)�mڊ���y>$Ւ�'��m���	藿�;���;?M��=�?�=k��������?��=�&����.?$��>�rp?�֫�e��>������A��>���.���z>sۜ?�z2>�ZN?��u?� e?x�+���y��6X���k>4P��+=Z>�І>�����.j�sp?�ŏ?�0�>��?\t>�Μ����pr�a5l?M;�?h;ľd⏽KVO>+��?`�1?vC3�0�c�7|���T�jK�����y��z�
�0>��?F� =��O?���?�r���:?��?�F��.G>��>�g��/ƾc�����ﾌcF���{�g�G�Q��q=�8�d��L�Uݾ &� 8{�����>���>{�K?=�v�?�F
?a?>��w?���>1��=��d���J��\��� H���>��ࡾ�Tt<gN.>�䱿Q�P�s����V��g�=��>�13��?a�e�`s7?��&�xN�>��>R��>)di�S���7�?]c�?�2]�x>�uB���~?�6Y�\��(��|=8��v+���E�ȶ=�Y�ҭ뿨s�0	?c�G���>��3������f�/O}��~:��/p��9X�6�f���C�������u�t?U�[�����(�' K=�*u��h���B���}?�2��
?�m���f���S>��A��j��ݩ��{-�4%U���)��3!�2�?�?�q��m;ʾ�>���?��H?�]Q��?r�M��Q��G�Z��?���>V�꿏!h?�K'?���}]��I?8Zr?kl��"���?�����J��׿
[l�7�3��#�v�F�>G�=�G�X�O���?]�u?V�����]?�7�?���?=ſ5k{?�q�?2�Y?����l��U�*�W>=�� �徍B���?v�{?*!�?f�>�=�?�@-?���?s0�?l󧿭�@���?o���3D?��$�K�"�?�󾤑�?[N.�q�žE�?w�:?8��>�/�~��3����ھb�\?�5"�
����"��W��{.��&�G���ku�=UvL��zG�,ǹ��X���u��|{>D��>���*f�B���#���j���6��飾�b�>:���ʾ�
?�x�>�ʉ�p�⾹R��.�s?K<�a��?�.��Z��?dx��Y�?H �?Nar=�|�������;�C�?Sf��l���5��9�?�7�3���J�1�w? ���S��^X���ϴ>�}f�b΁�S/����?]�����>��0���
?��_����>��=�`���k��<��D�ľV�?������>������RF���=�Rq�	�¿�s0���>��h�|������F\�>?���z�	�xs>q՚�L�}>�B��v�=���U?^?JS>.о����Q۟��p�>I��⯾F!�:�=Y# �L�D=���0�>���F���c�8����>WT����ʿ`&"����s�=9-"�����տ�{�>�޿����N��`�x`h�Q�Ԑ���}��K_,���<�(��6,��]?�;�����J5>�+�?k">�
?� @Nl���2'@��-�^����Pl�
8e��.�㾄��"�>ZX�h�%���ܿĮ-@���>Fg?�M�>�����͠?�D��^�?N����F��3;w�7�?O���;[���f�|}s?M�g�ǖ?yM|����?~!����Y?�Gy��]>ď��+?ܾbK��i�"�����=Η�����`���t6?B潿�\�>�����>[ϴ�=�R��S��`�>G�����?4�?�nq���>�i?�Sy?�E��+2�?G����?G=�;�(�>٤�>!�>X��>�V�=	�Ծ�L�>�����T�� �����>
�.?󺺿�]?�y>�f3�qȿ
S%?��M�"7ܾx_�1N�>̝>�=��<?��!>q��=��>�޼R��>�ý��|?D�?���?ܤ>�:F?���?g^`>�����gR>N�?C��f���_{��U?=Q"�w6�;1%@!p�R&?��u�5 ��Vv�L>՜Y�6��\u�j��������[��"M?��P�$i�[�/����i<95��{?i37�u�E?����jCu?Tb���T�>�ƙ��??�r��Cm���r�e+�>�Ⓙ�ĳ��`��8*J>�����Vc=�Y�9��>6��j�?b�)�"��?�ϋ���@��6�w�?ڥ�$�?#꫿8�¾�X¿2G}?�)ȿ�U�f�=d���q���>B����>ۡ˾8kJ?�b�8w?�<���i�<��1=��,����L%�>=~K�[���(J��	E� �>��*��7��	?��O?
n?�0G�?CZ�ݻ�>R�8�=��>ҧ�J�6?ﱦ��?�@�]o�]i"�չ�>�a�9�i�G�W�7��>1O�X�	�}�O˶?�'q��)O��W��VQ?�0�ی���=�:�?f���
?��)���X���.��f���?��O���?GE��4�?�ࣾa�����ͽT#�Rô�D8$<
�[�sK�>;����_T�Xjf���?qhr��#�r&"��ʪ?E�O���e��O�L�>B����ʨ;H��Bu�3�����ѹ�L�L����6��<e���4��/��d�>@���I�������<?���v,�E��PMV?ߪ�F*�������?�����W�ɾ�&C?�����T��ϔ?�s��<��>5^���*?2<�\G @z��?�si>q����3�kz/���z�VA?���1E*���>Wͫ=�c>��Z>�E
��2���n<�W�ZZ�=�P�C�x��!��t	�{.1�<��������3@���>�S��4��5a��۟>2�c��18?(�i�>�?Ä���i�?T1�=�4?��>�W�>�����i�>V����?|������iG?�ľ�M�=��+?[x�?7�>M�F@D�?��0@ጀ?�:�?\�=Ht2��=n_?�|C?�=����;@K��>A�?�*����.c�>���ࢰ��m����+��K��j��	��U�r>l�οRa�.C�=����Y�(�)���_�e���(����1������5l=$�R�mU�k��]����(?C!����3>ԝ?�k?�?��v?T����`<?��>��5D��$�z.�y�����<�N�� �����ͽ��)�|C��K9	���վ ��HdB>�E޾kQ=���Ծ�^վE��=��?$6޾]E�=oǾDj���0����{���W��0���q`��n�ʘ��? g��p>>�,��?���>�t?�þ"g���*��L����a��#2���.�H^6����w�
�Tj�?&˽��v?69?�ʲ�+y?<+��3M@�����?�U��H�P@�q?��s?Qf̽s�V��� �m�?e���=7fo=�x:@�OC?s�
?���>�JU?կ?���?��I���뾘�ɾ絋>���=���He8>���<��a>�����	��e�eGw�X�]�]2���d�<h@���
��t��=���1���/����Z���q��|/��4Z�>����ܪ>�z��5l?����}��͐?W��?&?"?nţ�4/�?xl�J��?<-����@�'��򿓷�>a/@`�(?I��>�!��OƲ?*G?�N�?�??..�?1_I���X?��>*[?��m>��>ݛ�?��4@�u?�0�?��|?���=�1p�!�Ҿ,s�?=ZK>U?a�?g_?���?�?�?�˸���>]r��|���X~���Ѿ7�5>���������k��Q�>�D�>��>��=��=�-�>E|���u�����I���<��G��e�
�7��> ��>�V�=��F=-彣 ?몗?�E�鼧=��&�*�羬�?V=������!&??��>tG��0��H����>�!�(�!�b�a����vjL�'����2>�Ά�����ܥ�^�Z��O����1��:�>NY\�ļo?@���|�?��	��7T? ������?9N����,=�3?4`���;�Nr�=Z?^UK�X��=~��@]=lQ���:���]���=��i'���w��'>����=3?�E�?7�I�����.��3����P�qW�>�?��W3?�;E�?s=�ca����=H�����L�^��ڋ��sp?���7�ҽ뺿��T?C���r&>�=�K�ɾ�����뉽��Z>
��<{�?�>Ml��3NC�sǦ���H�n�Y��WS���>B0R��U�Ⱦp?sR4��Lܾ�<@����@-Կ� ��߿In? v>{�>��?�4,?E �ͫ\�A�S�%e�?�UE>5�R?V��/�?:�??�%@$g�>�i@���?+@��?��M@�[�?���?��E?g�@>���?��@���>�*;>j��4�?H2;�۞��Y�v�VX?沌?��G=��h��?���?��>s���
�>�
@u��>0\����޽4`��QpK>L�&��y�Vp���?���
+�?��d�W�?Y�M��=�?W�?C�>�?.���Ci??�e�?��-��b���Q��zq�?,L^�I1������-?<� >(ϔ���U�Z�Y[ľԎ�B����?h��	��>꿯�^�����*@��$���H���=ɧP�Ȣ;?0��U/���@��T���QY_��v��U֔��ak�X/�}��ِ/��z?����
?^7	��7?�4�by$��A�>~���?e�U���>g�9��3l�A�V��T����3��ȉ>?��ߗ��q���	�$�?�D�>��<�NV=c>v�!>-�>�2 ��'���Q�L��>�!��KI#>�xR�z?r�<�>IL�j8ٽHN�>\ݾ��3��(�W�>/�|�ǡ�>��Y�W�)?rGQ����>{�v�T�.?���>D��"7\��v4?�+����l-�?��տc��?��U��E ?�2��@�?�I���_e?+����о��Ǿ%�=��y>5m@~r�?oG�?�]��&޾�ɑ�U�?h��Ȳo��a��@�Ԝ�Wl|�u���1��?�p��p��>�b���.?kk���hоL���1�>ӟ�Ԫ-�(\���b���瑿	ܚ��w��S#u��B�Kt׾��������Ǳ��X�=^p����m�v��B��yU���
?Q�xu�����>�i}�]�����⟿Ȁa�u�`��\k�F⍽?l=�M����l�=��>���> ל?��b��,?�T�����QX�2`�>��w� !���ǲ���^>E����ſE����S�qzm��
����Y=��W>�Lc��ԏ?�����9@�b�O98@�H��an�?=�x�z	@�ѵ���8>y���f��?߻��xd����O�>�%?���+����U����_-?��Q>�i�v%?.Ev>��h?�?�??�#-?��g=X��=3Bһ��>�¾$rF��ϼ�2J�vƋ�PzD�;�M>U����E2����>a|?�<*�|)þn�p?�Z�?�k�?����x>��k?9R-@�^>��@�t|?��@��a>�FG>V
������ҁ��#:弔�3>-ǵ?5jP<;^`?y�N=%�+?�9>�r>i�>NH?}�A�sS�>���?QfƿQ��%��
�t?8(^���J���Ӿy�=P�:�_��?�
�?�+�����������>�1��Xݿ�B�J��2�>�@g�!���=7N,�I��?��L��>��?sb@l�1���@	K�>��?�.��*~��6:�0`^��O�����[��8¾I�P����?������V�I8��y�?nt_�$�6��X<�w��?5QH�7��BL�h;ľ�9�L;?v>@�J@v��+&,��,ￎ�Y��A���'���aֿ�ܿ�V��F]@U&��+A���B��1�>1%�?��־����p	�?Lp����?�u���|h?�;�?���?�#?���>�U4@6� @�:@[Ҙ?Tz@�}Y@``@Ji-�$R0�G!�>Jf���8?��&�!! >&+@b��>4h~�}G�?��@��+Z��گ���L�?r氾`���^>w6�;���>%�L���@���Wσ��*d�����&�4�X�����8�'������� ���?꺿j�@��?"�����?����,�A��#-�}�?#ם�Jo�|�4��>[>��&�>[��r���I���悿��h>�ȿ@����LF�9�@�m�sue>6#?�O�@f�%��OY?�nM�<��?�����u^������,��t��S,Z�֗������Ɛ��t��d���U������w#@\���=�۾3� ?�R���R?�׾��?���%���-!�@����ҽA��x���ߙ��W=y?T�Z����D��< т?�*��j,K?QI4>GC�?RX���
z?E��>�"-@�ѝ�>�?�,?�1�>O��? z�>Ŋ�?��;�~��?��>��]? �>�O�?L��?ߤT?�q�?��?���?A��� @U9=?]�@,�8�gJ�?
Q@q��>R�� /?Ÿξ���<��os���?a�Y�2�n�æտZ3ܿ����Pq�>M��z.�{����-Y>њ�?���"?}4��};@�i�Vy�,����M@JF��58��
�f�O6�?��A?ד��sW�~�?+����|��O��՗Y>q(�l��>YkF��С>�<���?���qS����=7��?�C�����(��,+�?�.���7��!9��
?"����;��I;�o���+����=&J��Ǫ��I$����zN>�f>U��'#[��ٟ>�|����,�//�=���?���>aR�>;@�^;=ya�>��뿜{o?�*�=c�ܾ���L/�B��>mb��+{�<A��P��ޫ���.>�:�!�ҟ!�?Ua>3�Y�A����q�>n�>�o�?��>�Ԣ���?�H�?B�>�G�/C�?m[�?����ѿ��>�U�2`�i�?�.����ֽ���=��e��+?}��>�b�>j��>na���7���E�=%;I��<�޾XP����0�~�#�7��}:�>Ԑ.�9��l4�ƀ�kӾ*���侜)�N���h����C�>�.۾Ui"?x�1��s?X��>Q.��?��?Hb�?J�?��@RP,@K<@]R�?nr@�@��?�q���"@�[�>���>ɑ�k���.��ͦ>��?&��?�N��Q>��B������B�=���=/��>}�>қ*�T]>>Eu>�ܾ҇v�/(;?i�	?�Y�>HC?�B>i⵾k�?��f=�~Ⱦd�=O�&��Ծ��?�18��tU?Cċ��~?ajb�WU�?z,�)�>=�1L?��O�>Y!���y>>�����1�_ U����<���=��=J��~b�f紾u�P>���)r�>�0���R>H?��]�G@�1�>��7=^���M��p_�.���𙽵E�$/��H^�Ɏػ�G�<�	�;�'�ͬ��	�>�L)>ǒ��7���*��V̻O��=�3,=���V>Ӿ�������f�ɽEo?�з>�ٱ�s��=���>J�Y?����t�����=n�F=�1������9u*��h���c>����W��>��پ�?�&��Zz=h_	��\T?k�Ǿ�W�>e遾6u�?HP�>4`���'��#6?��P����4a�o��>94����n?.�[��(�>e@������=��C���=�ݾ�K|�A!G?=�g?���?)R��Nӽ>˩?l+@g����[?��>>
?�'�%?䮳�[B���p���̲?C+�>^|o>��=�RS?W�y�N>�1Y��:��U�����=��q?,�C�h>V��>(��?m��?�<>h�b?_ G?!��?�>/�L>�Λ��g��Ң>�������s>��?�;�[:?�s�#'?�q�?E��?s��£��\����v?���7u�\4>��&?u����L�nD�<4$7>�d:�������5����|5�0�ܾc���j����+�
������:a<Y�a��f�L/���Ӿ��?Ҡ��P?����eK������i��j^�����y$O���I<��g>�����y��u>O�g�Io� y�?�~��&���)6A�x�E?w�?�>K ?��?M��?#th?��j?�2�+T������c>��R>��	*�~[�>�J?«�>�!�?b'?
>?�}�=u�>�j��7]�ϹC���	?����:�8P���->k���<��_�>žz�^�CK����d�,V���D���ݽ�j�ӳ��D�_I�=U��>jݾ��O�����D@��UgW�?��]�G@�M=^�?vvX�	~?�Qx�S�?EM˿�-p?�ݱ��l7?�.
?5?�^k>��V���ƽ�t�?�.)�=�>BJ�?l�?�'��Hr?5�e=��?r���.�?Y揿gZ?�`��Q8?ɇ׿��Z?WZ2��-?�͚�q�Y�1W��4N׽7�-�1�"�U�[��Ц>��ܿѥ��9/���.?z轿o7�?��^3�?Jz��T�?�Yp�� ?��Y���]?�
?~ט�VfN��Q�� �;im?�����T?�O}�R�o?������?4@�?S[<�e��H���Ik��>�8��@%��^���(�>��V�F��m�k��̾�Y|���f���S�;�.��$��DR=M���0�� �����<%���z��~z)�,h3?�؎�	�>1�����?{���V���G��?*����D�ׂ��]��>0F���L�L�Ծ�p�>�
������>f�Ӿ�п�ۛ���@�hQ���?Km~��F�?�ы��'@�;@�>c=�7��H�=lv���>�J�68￀���|�>�b�C9�HX���$�gf�t?�����?r}�>;w?�m9��Š>�?�~�k?��=������)�7Q:�����1@���2��U��Z|.�����9Z���F?�*.�e���-#����>�9�v,�L�8����>l�\��� ��n�ei]�Jj���@��k�??������?�]��}}�?�������>?���  '�Ѳ�>3׻����\a�(������u�?�ن��r>77���?����.�N>W.���ڤ=��Ŀb�o?��s�V�?����Qpa?\Md�dي?}����?�%�l#n�뀺��?5|ؾ�8��mi�?&�u��"\��EQ��)�>1 ��ؖ��(�>���>�,>w6�;9�'?e��\�����=�S�i�?9fF����?�_���@!�����r�l�����H�=�a��,(���X@@t�>;��?7V?M�q��ǽ:Ⱦf?�X]�[��>�J�	.�=񒿀�F��]��A��>/�x�#?���8�=�?�/[���=>媽��>�ł�'�G�lK��W=���?e�`�b� ?*�7���?Q
�� "?�Dg���?��]�G@*��?ꑀ�i@�b%@5�1?)�?L��?�`|?�qg?F�a?D>���R�?�(�?�vR@E��@���?�Ǌ?pD|�g[?a2(?��H?��[�V�>��?�Q@L�K�j�1@���?��@twd��yJ?ΔN?�E�?�Ⱦ�??���>�?q�q�#�Q=j��Cv?�`�7�U��t��qm�IC��N-��<�����љ��v�g�՚��`����(�^��sS�>�^�?��m���'?n�u=#k�>t����̽�0b����xPl�#����������4?��L��r��;�O?��;��־V<9�=9)����>W�a?�+��F~���S��T�=�
��.�C>�� ��(i�SDD� �?�R�����*6 ��1�?A���?>&`��#?4�7�V>�C,<^�j>��,�>'���6�����V>��&�}���`'�T�>�V+��H"@6� �iD�"qK��4��D��ޣ��&c�?7�>��7�T���"��x�1#�>�4C��ga��u����� Ep?�n?��h>7$�j�>��?��>z�O�K޼���?���0Gr�p_��V?G6�?��=>��?l5y�9�=˨�f�B�
�Y��v8�%x������/½^����>��>�������>0Y	�]v�������Z�>k�n>z:ȾT������q����L?ʔG=��վ�N����	?�j^��su>;e4��]��>]���=˪�?N��߂j�� ����ᾌA�>�hJ���?$ݎ�[ܮ�G ��)���q�������@����Tl���.9�Ì����?d�����&@U�C�Ts@���>��@t��� 0�?eo���2?��l�"c���U��u�����i����<�����?�<���=� ����?V�ſ
Q@f��86�?Z�C?�??�����P5����\�?kk�%?���6{��ž>sN�?� �>׾]�J���N޽K!?�*�?=A4���>Y!���ȓ����=U)�?R�?~�4?u�?ϒ'@B�?:�?�Ĵ?ȉ�>��>d�@a�?�u@���?tמ?�+�?.!�?V!.��2�F���o�>�d׾ࢾ>2�!?��K�eq?9��>���>��-�W<1?�h�>��>/��>�\�� Q��	|��g��P���o��SL�=���Pž�u1?��5?����}32��t:�?�?��վ�Zw?�g���f�1y�;��?���yd���.�D�?�`����{L�mC?��3��Qj�����i�����?�3�4��u��Ea�d��[��,�C�e�k����S���Y�sl?����뼿�m���]�?󮤾ݤF��s�ꢄ���侑g?L���wF@l��7X�?��8����>�H��G�?@�>ҕ�> �TAU�+��i?���w���*@m�U�H�@yC�i΃?_Q1��+.?�����b�?��>w�?��a�P�@_��>�p?:�>���>���?u�@��o?5`�?#�>	-�?=}6���@3�g����?�O���8�?���ή?�ao?�j�=1���A�=M�o?�/"?���/SN���H?ȜҾR��>��
?wG�=�����Ᵹ_��8�;�Nּ8���5?P�?i��>�>�A>K�>���>�������?O�ھ+��>�����U��\���5��A@��'��0�����?S?WJ�%�j>����ą��.���@����fU?&:���:?EžV[��v���@z�*�ؿ{lp>=F�?��4�6��e�N>%y�>ƮG��hʿ�Z���
?�9��1��e�U��rb���?�g�m�d>)F�k	�>����u?��v?ܻ�>m�t��n���3�Y>�2_����b�*�>��u��{?.b��^��v�B��T�?�>���x���׽"����{���w���ν"�s�{T׾� ���b���*���-��q�0�������?*������y���o�>�����꾤���5?)0>��{=.�>���>/�>����P���r��E���C)�����n��M>���ϼl�پ��о����<�O��>������)ľL�#?Y�.���6=�Q�<l��{��=�ٛ���f���F�{8˼��OU��rҾ<M����>�q>��-��ر�^Pս�*��u靾�"�� �8oc�Љ�*�� ��a0e�x䨾����-!���<����h�T�#�9>�w��� ���u�U��?�m���>���c��?󕑿�(�?ڪ���@���Ҁ��ȳ>�ɖ�G�������b�:>|�?��?ߘ���#>�5��h��?.tg��*?�c`����>/�Ͼ*0�?@R=�D4��y�7�T��?�td����>\ƾ��r?/�= ?Y�F?�L�?�8>cu�?�ƈ?T�?ARA>�!>�?܎�?ۢ?�D@u�(@>�@`��?�h$@ꢄ�<k�?�Տ�!�>F}<?�)���v��b0�q����h��|l��b���{���T�;=?\|8>��6�ؾ��=����=�Jwv��`\�W?{w��>�?���8n�?e�=^�?+�(q�Ր� �?
k�=h�@?�Ǟ����>���*��>�@�r��?��}>3i�?�	�P��<�!~���ݾ�R�7x�J֕��We?�8Q�*��8-�1���4�	��}�?��?����C�D�=�?�t�����ې��v�<P1��&������½	�潾�
>|j�=�F�y�>V��=*���,����ڿ�fa����>���k�?�:��Ͼt��Dc�?
R]?\L>����e�?w�����>t��^�?OS'?�|@>�S(>��D�)���|��bƾVd�������l.�U�B�*\��߁��%�;~-r������qV�>�V<w6�;^Yj?�Ӂ��IY�?3��BȾ���{���_[�Й:�כ��3���TE��'q�=-ž�x��Ё�����>=�v���!?�}M��nԿ1w��]@ʁ������Z�/;5?&��z��ʡ���n?o�B�3D>��C��r�?8���ԟ?04����?ϼY�� ž,M�r,?O��ȅ�:r�rr5?Y��ꗻ>mk����)?��ikb>}#��q~�K�9��Λ������3�?sˬ��P?�5���@�?��󿳧	@D�ѿ��?i�پ@Ѿ`0�?�������W�=kF��9�*@��?�^@q��Uׄ? �J>Jk)@2��=BO~?�#>�r`?�N?D��>�Ew��l��g?�ә?ٹ�&����@�-�?��?�?�?���?�M��Ε����ez�>.H��ȑ�>��$�?U�>zW�>�H^=��?���?P=����>|���5����>d���fc��d�>C��=.G>?��>3��=?Q�>���>�o ?����ćA>C�>�?r6�=�_����=����Mb:3B[����=��?=���`U����=ݖ\?����c���z>=>�=����j�%I?XFG?���>��A>�|���U�>�} ���'?�Ģ�E�?0�����>p�
�a�"/�>1˽f4����=�f�>M�?�
?�{H?[ܥ�뤾�����ᾩmt��ѳ<��������w��\@Ⱦ^%���L[>�ƌ��㋾j�^��>@(�l#�>%�����bi2���ӿ��7�X��w�Ԧ(�����F3�?��6�Zߙ>�S>W��?5�>7Ύ?c��>��?��Ͼ�l>2o��O����j�z�����o���pˡ�T�?tko��-�����?{����O���>�?�^���U���;�ho?���[0�<�E�>^w?���>'@4G�>��?&�7>w'P>}��?����l��*���\`�%�@?r۾D�?�ɻt��?���.>��l?�h?���3\>�J�>���A �V6�?�I]�Y�?5�)���q>>��>�C?��'?u�?F��>Я5?�����>��˿9�?�Ρ�?�?HG��f�??>�>s����O?�XZ?�`�?�U��սܺ8�.A!?��A��>;?�fM���?�E��Gvv?T��=�W>˾)>���=e��j־��?Ŀ�?�8T�R��x&����?s ,���4��I�*�a?���ꉿa%$�u�>Mޏ�������9���ݽ�6k�����<?�4�r�'`W�b
��IX;�z��=|K)��T�FXG�6P��ϵ'��\��E�4�q��+/��f&=�+l�)l���U�X�B��}w��� ��4�?��>�c>�w�?��տ�`N@f�οg,�@��˿�@˄��ˋ��dR����>�?p4�>	�+��Р@Q��?�i@���?���@wy�>��@3,�=��@@�H=��A@�M��"j�@d?9?�G�@\��@Pj�=p�@XO����@�0��\&@���?d�o@망�Lt�?�(>S�?�����<��?�^?��S�t��>P�r?$�==Lt�Z�&>w6�;\����޻>i���A��>	�������V����f^�\]k�����!U>�Xm>Eb�`3��Ca�������>��$�LC�>eE��l���̏)���Q�U�W���V���/��
T꾑���;�é�>�*�L3�<D<�)?����v���(>�u읾Y�-KI� �u���/4��݈?;�:�܃?�v�>�@?����-y=�5z=ݫ>��}�;�ɾ9�)>�U���
?lA��6���>P��P�?�~�=�s?���>U�n?P4�=���>;9�>��<:0��A"a>�����"������n��]=>]�*?���h�=8�����>_R=�,ƾ|�y��Ӿ��۽J�;������N�>�ξ�x>�m��4�%��@��Gz�=$�?7:Ծ_'�>9h0?�tC?J�� �>�(�?{��?�ľr�>�V>��?���ƿI���>�M��
?X+���&�<hƾ
6���
v?G�b�"�?�V� ��?�mX��|������Ӓ5<�DƾVd�����Gȸ>�\ʾ&{?������ڄ?�50�/�J�e����?J� ��Û��kT��!&?�GR��q>��8�	��؍��rFQ�)��wS���f�U�NL��I1��q����!��k����S>B?x���u��˽M�>.�.��{��!����޽��=�|���?��S?橾����ƨ�>��[>"ls?C��>�3?�|	?#�+�&ɘ��k�<��Q�t>�(����>��޾�A���׼�k?�(*�F�S�5�9��,�>».��̅��<$� �>iB�>�$��$�Ծ�E2�q��ΞI��p���@���='�����>��d�U�����@���c�HI�)�/��e�=$��嫗���Ǿ@܊��m5�P.���� =������� �|��H5�?�i�=;(G?��^�b*<?/,��3�>[zh�'e�?�{��z��m?0�?;���?�d�	�u\c?8��?7�&�����JĿ�Op?��a�n���v��.�>*�/��z�>��	�[��>R"����8>��H��h?��Ľ�>LN�>�>T�=�\�>$�?�>/� �Oj�?Ӑ�q��?�+ɾ~V�>�_K=��?�&��~>���K"���
?�*������.�z������eL?>�|��,�?"P��uS~?-���󩽤v���~=_�B�hC�=!Ռ>�c[?0�g��!�������?��_���o>"��:�?����r�E��ܾ��>�i3�:�(�BE�����Ǩ#���ԾLa�^|��8��^��$�?�Jȇ�3]��i
�pe��﷿����,Po���n��eп�m7�<k�=�-h��d��I m����>�`p�Io��+��~B,=�>?��3�^m�>-r�>�K$?�5�py�>ſP�Ǐ�=K^�=���=��.>����w?�D�?��C����O��Qg?4�;aW���׾m<W<��=��!>E�?�6�?>�?K��<���>PɄ������k0��ߔ�M�g=^�f�>v=��(�I�A�Ӿ�G/�I�R>��ľ~��%|��X�'�P����4��?$������Mb��� ���E?��$���?W��-|(�C>�^���?=�8���0?ti���i���� >g��>��?ѻ�?�h��᠈?��?�>�?v
Ŀz
>����n	?2� ��\?뎕?5���̿��=�2X?��?�������>L!��n&��WѾ�޾��pM/�� >+<��ܑ�1!�.f��K2.���@�_(���c��f;�w!k� �!���.?��>��>�u>b� ?g���Dh?P(?>/��>�>[9>z�>L�h>�)�>���>>�U>������(>�[��E����a>p^M�Y�>���>e��y>f�4>r���>�6��!�A>����J=L���7��eƞ���>e_�����>��>���>iN4?�h?6�ӻ��>o��=	�^>dH�>��>	�>.D?dT���G?P[�P�>�Y��E0?3~?��H$?�U�G%�=!8��5>�H�>`�?ON�>v��hĂ�s��=�z3���?��?�?�> dྐ���� @�f?]ʋ>�RK��>�Q�I�>��:?�U2?vZ+��o�>Qז>���?��KQ�?�"�L��>a�B�ψu?��˾��	>���>Ȣ�?��d=�A>�P>���>d���04>�=5C�>�ܒ�i�<>�>b�T=�d�3l�=��>��l������ob�sS�>C9����>��T?�Uy?�>��@ڟ�?���>0�=?;�?!�M�e�7�ڴ�?���?Pw���%�)�>"�"������?Re>���>B�ݫ�>]��>J9���M�±�?X�?�@���?&V1@�?Ӌ�?�>CO�=��v�Э?G��=H�?<�^>��?(��?\�?�Q>�G
?���>�w�����k@��wL?׋�����q��*U?:R�1��?�y�	��?0�>gd���A?�I��pU\?^ۇ���r?�ԃ�`���M�$�g�6>:{>�E{�<���*%?R᏿����O��!S�?�����>w���C�1�M�I�&�\d�MZ,?�T��?C?�$b�^S� �>"s�>� �X#�>�U྘��?�;�\���)��"8&?:�Ӽ3?����
Ր?ڥ�����Z$�>�L�?���H��?*�˽6�?/���� �
�=<,���e�#$U=����w�w�y�[�>�CĿ��@���I��!�����V�>(?�h�=����?;��?ʆ����?�����K�;��?����aW@l\��?d(R�;�D?����7�2?1(��+��������K#���<����>�����8�=�`/�L쏽���=&���rC������)��{5�/�|�x�D�ҷ���m���U��	/?�����홾!�8�:y?�{����?��y�ʄ_?��d�a?�!?�a>���F��>x�W�ĵ`?oŁ�3V��S���\-�?T_Z�`﷾ ��t��?{����e��MW�� �?z���D��*��B]�=�y��?�N�z�����\�j�[@���Q��xB�e���K��>)�\�4=��Vnc�� ?b�~��
|�E�,���>M�L���J�c�?�9W?����
?�-L?ǡ������j�w#g�-Ƽ��$��{��4��bt��U�>j��>mm4����}�>����A>���Lg?�Z�?���>��?Gm���B��I�)�@i�Z�{2U�`z���&?��s����c�7��U�?K�v �>�s�ǔ�?E-�,�	@�Z� .E?I)�^��?�!>[h<?��>��5@@^0��ի�Q��!&@�yT�(Ŀ��+�1��?/���1w�?��?��a?��?2��?:�P?u��rN�?,a�?\�?)�?��@vb@q<��K!��������M������?���>#�0?�n7> �%?�����^�?�>>J�=?�?c�"��?�@���>�@�"@ų@���@G��@�ą@]q@��f@�^?@?r2����ݾ'w��s��ͿX;Q>��?�1u=t�k>n�?}N�?�Y�P��[D��
?Y��j�?n��,w,��]x>���]9f?����?Ze���5�/��/�/��e�r���M�l?�>kȚ�Y�ӽ� y�K
a?�D�<�F��F����"?5�>����ݞ� І�+X?�[����ƾƉ��uMS��>�N����������Zr�>8W��6R�l�ľ42��� �������h��8>�X�xԅ�����n��>vyϾt��>�ֽ:�?�9��4`���V}���H?&�޿����Я��7
?��}>�?�g�=�I?En�����y"��5Ó�E�z�aҤ�$�����r?d�F���>�M�?g��7�>��ƾ���>yU7�q�D?�H?��5?R"�>J� =��O=�f�>d)�?��;��p���������8>>���>  ؾ��	?���Q�S>�\O�@t?F[��e>�+<=#ó?�;�?�3U>�I?ק�?,��?sS�>(��L�1>�ڝ�NE���^?�]J���8?�P��~A?��q�L�?9�?q�*>GrL�v�<���>��?&b�����e�	�?Ŷ�����y�k���<c4���?�L��e�	z�����f�ᾷ���9Ծ(���z1�vΪ�Jg����v, �d�V��3>�c<>0)��YO�%����?�L>5P��'�>�a�?�vz>��d>w7�=n��?��%?��v?�c�5c_��o����!��?��?H9%?�V�?��?z1)?��?~�?<�ɽ�jg�KkR�N��� þ����5/�	8�>�e�> ��>�zQ�<�?��<n�>-86?=��>YR�gl���%?�;{=s�J�^a=3�ξ6�����Q��>�Z��W#�Z�!�쑤>3&�=q�> K4��?/"E���	�����<� ��ԙ�<4iվ������M?b���U��Yn��轚���J�� ��8N��3��پ��'�z��np?�ur?B �վ�̱�?�3���g��B���6?X��5/�]��y�?�<e�t�~�q婿	��=~����D>餝�c�)>����^��?�Ú��榾I�u�1��>mYc���a8�"� ��Z������(�ր�X�6�́�=��Z�7~m�0�`��Y>>�c�q8��i=�bN�>��M��
?V�׿�(������������@��ɾ��@���Ǐ!@ra�v!@��@	�8>����ƫ=�"���i?m����&¿��T���?U�6s��b=a��[�?~��=�{������pg�Q�>J0�P����4��i�!���& b���j�D�L��o�>�;��|S���;��N?�7)���4���j�?����\pr�����Ap?��&��⢿���
2?z"P���v?ŋ�?4f��:�<��rپU�k>(��>$>V�<2	��w⽖��>eڑ?���?M�<��$�Z`�;I���C��>茂>�s�=���>㿒[E>��?�;���܇���0����?��Ͼ�_ƿ�᳾7��?ڶ�)P2��\���e?�Ԕ<%uҽ�l�Z��>2�&��+�?��s��޾�=5�;�@$�m��jƿ�����@?`r�T
��p�	� @˜�� �ɿ�˾h;ľ�@=<)�>�s�n|����=�EW?\����9�����cO��h\?�,_?����E9��ۀ�.���]e��m<����
=>ێ>�3�3R@BXD?2.?���?��?�~a>�,�Ց�?�8m���>���>^�q?��?$T?��@W�<?o��2)>p��>��>�jὰ�p>��˿�&?�ԭ�'/>w}�?f��?�s��Cc?K޿��="�Ҽ�I�>w6�;&U�?G�����?��J�3��K��ױ-��[`�`�˾�:���n��xw��o̔?|�?Y]��f@>�J�=6p5���'?X�`���>;�k���4@K�w�'�	�`�J��@��O�vC�y�4���?�6��k*��oA��?�b�`��>�������t����>I�"�����@$��?$7�6��Y�P��?�[�Y���e����1?U�������]�R��U�&��?���b�A?\�G�"�_>��>�M?�>�z?-�??Ȑ�����N	}?M`�=��E��;?"?������x�/����?,��{��>�3�=2��?��b>�T{>�}��P8���F�~rF?tz��4b�?Z�νv�G?E� �X�����D��??0��wؾrb��������ȿ��C���>��ž�7�Zc�=q����뾪�d�a�5?�ˑ>��μ4`��564��	?A;���B<���?���C��?�Y>�k�?�uh>D�?��	?k��>����༤.s�4;> )>����� =g�Ԧ�?�*�>6�%�%�7��k�?$蓾�up���1�uQ>�r)=S��>��$�.>�&>x������Ɲ&> 0������}r�r_������o9>؍��f���L,��Sɽ46��ڽ��@��?C?�O?�@�u?�U��y��*�?��??��>Wrt?�����τ?��?4�?�{*?�np>�A�>�,c<�-@?���>�~d>O�?9��>�\��&K���*?.`����ھ�8?Zbw?u��@���>c4^@T��X� @1�4���)>��?jC��{��?nH?[�@o��>��V?�P$?,D޾탂?i��>�т?<h9���p<tީ�G@_�
�eKy?c݇?���?�KN��$?*A?����h;ľϦ6?�5�=���?f}?(኿i��𫻾��=�de�D�E<A*�����!�'����?R�>�gz>�盾���>^�?�����%������_?��>k�`>ly�?yģ?Zp@$�^?`_�? ]�?�89?s��>H9�w��<����!=�8����7���]��`���4s?�A��A�;?�>�.�?-#>m�Y<�s����>SJz?P��B��?���?�̉?�U�#��=��.����j�6���4���N����Ƅ=7+?����<B/!=
$�=�[ľ��U�J�?�� �P>���t0�?���<2㥿Te��N�>(v>��H3;�IJ?Sh���o���`	�w�@@��?"g�>�Ծ���?V/?�ɵ�W�D&?`��E���G�-������J��?uu?��-�:�A�	�b�������\������ూ>����'=�U���>��?�m ?x~�>�տ�n�=~쾿X�ݽ�r¿%w
<7
��_~��CI? �?�5�n:C��\~�5�½2�?�Z�?��D��@���o?�	�=��:�\��<�?q]��� >�@�?.>#��z�>B���#F?��ľ%ڍ> ��>}؈=��>e�C?
��?(�?Q��>`��?�e�?���?�-W���@�0@�P?�Fy��8,?6�+?N�C?�޿��>�U�K�[���?���?ܸ�!�ﾏLZ�4�?��&�?��PiɼgA��?��&*<�>�8��or@��?x{T���G?=��M9�?U"��䖿_�^�eԁ?���i�|����,�F?[������A��S��?0���\V=܁��KZ=�Ў�Le����V>u�M���b�ܾo?�C-��8G�q���q�r��K۾�_P� u?Z9�����ʻ+�5R?�4���U��Ƅ?"e���1���>�p?Pf�>7 �?E��?Y�?f� ?�fֽf짽?,?���=<:%�g�&>�)����>�p����f�?sF�?P����>h>ϒ�<PHI�P�?�v�?�P?�*���S�2
Y?�$u?΃�R�V3?�i�>!A=�"8��l�> �D��}
�Z�>>���7`�"��my=*��|�,�坕�W��>u�?_��(_�>WPT?�?�� ������?�h�?!��?���̠�>#,1�%��=qV����?�֡�P�����Ļ��?=�>��$�Z�{f_��t�>���=�G���x?��)���?��?ߧ�>�D�>}u�?Zs?�{k?>�#���>��5?�H�?�U#?��?�@,$m@W!�??�Q@"Ϳ?.,@�?#�H�?�{����@!}��H7?61��L��<b�f�b��?Dd�=h�|>�8Ǿ��sS�>�'?�9�>Zþ�D�?'�׾KD @�|��a�?o����$@k.������
Ͼ}_�QV�>�!<>cA���Z�@��;�{@�y<
;Y�J�ھҜ=��m�?��7>[�6�0��=m1?ݱ��J̝�D&��e=��������E�H�X`o�C�S>#j��;�>f꠿�?W?���Yʾ���\�徺�R-�����`������M�/��� >�m]?�HO?��v?�`y�_��?t�����?
����(�>BB���u�?S�?���w?����2=��r�3=��'?�
�qٿU�����?��J?&�?kZ���s��a�c�H�������>�@?⌎?C���v���\�?�Q@�����N�\�?�5�@�(?��?a�@y��@�@/��?�6v?�o�@u�~?1�@���5�H@��?{3�?﫰�a�=]1�?�)@u�ӿ삾��H?��?3��� 88?Xª�H�n���q����"��4�S�#���n��Z�>��X?�����۾���O��?gG�<�	�"�f���@EA��G���"� u�?Ǆ����=3I���?K�B3 @���#?}���4?o.���>�����9?fH����(���L����=L�ǾцK>
p���?�`*�̖�=&�?���?��[�1�U��]Ҿ�� ���m�	��?��|��w�?[�����$@%%��g�?O�����4@{b��b���>^��>�f��g�L�[[���
@����K?-Y?��>
ڻ�>�����G@r�&�X���2BU?�с?a�$���>�H=�S��?cz��.�>�:쾾xl?��q=w�<���}>KO`���?�������?s5>̜�?�@� �?U��?�6@s��@Ժ�?U9@.�?�)@�U�����ˡR@��?K<E?}�^�p���t�z�?U�*��W�>�䛿4��$'�x�@�C�?�Q>�~��ҽ���>Q2�?�kA����>�?>��?�F��ɠ/���=D[�>�T˿��P?�[�.��?��M�N��?���?��@C=@�B@0�\@-�l@�O}@�a2@MB�?b��?��6@NQ�?����zX@LÝ��2�@*�"����?#�#@�^%@��&�v�?sS�>V@	��fZ5�BB�Z>>?�"��G1>!h����>+�s���?��?��?�]���Ҿ3�Z���>M��=&��)���h��:پ1?ౄ����?�Q���	¿�b"�)HL��䝿h�c?x���)?�����#�>�N#��?�?���.pW�8�_�2���u>�l?����9xL�������!��R�g�;�D����>dO0�W���=�?�u/?;A�=����:N��)?_�B��)>�?-ؠ?^�0??P?��?��?�O?�R?^z��Zr��M?�=?�䚽>?J�@��?�r�>�۽`#����
?�d_>��
?�� ���'?�����>C]��$�?�T<��f?:�ſ��>,N��k�>��t���?3z��f
�>�9?�hC>>0��Rv�>���=�ݑ?]n�����?�g#?Q��?��R��=Y��<��?�U��TT>`<��!@�X���4?Ry۾'֯>^j��1/?G-W�ދ�>z �>�D���@���>��@� @��7�����!��=\�>)���z��cO�
�i�����?�*�s��>��	�>�'���b�?���g���-��:0��f����; u���S?��_Ŀ�;�ݚT�<���fO�$Ӣ�
� @o����J�>�UD��� @�ܭ��Yn�{�I?ꢄ�kM;?00u����>P���?������?-���ܝ?r�^�伞ꔻ�w�>a�>�'���i��&C?ɥ��<��:��=�?�Ɓ��������%��=�/���s�����Y��=/�0� ж�z�s�����>}��T
>�xa�x����<��x�s?.9�[�?ͨ	�K-@�J(�?��?N+k�&�&@�vT�5�?������?�33��C��n~�m�b?��I��Λ���3�/�?bsҿ�b�<��?�N�?&kg>�t#@v��>���?�1H?T�K?��=w$���*�a��sh��y�?�2�.�?Y0�;�)?�� �"��>`9�ch?#�h��V?j���:��?�b� )>'ߑ�C�4?����=�񺾹!?�Ė�$��<�c3��(2>��q>��T��Ǿ��^?���>��>��d='?rC�>�B?�2S�nE�?��$? -�?�� �]*���@��Ծs�?����q}?f��5?�����Yr?׫Ӿ8�ʾ,�1�	�>��.=v<���U��׋?�?Ѻ�?G�ؿÃC@~��>0�?ģ鿰U#@L>��@�;��(��?����0�?ܣ�$�@����d@w7�?6@���?�w�@�A@�@=?��@!�@�XA@'�G�%�?K|��G�1@��>��/@�j�?,@b���Zt@w6�;���?b�¿%�?B�[����?nG�">(?�+���t?�S�߄?�]�?��	�J�?�:?�~���?�CP�'V�&]h�a)c��ѝ��(C���>G^g�+�=�=��\�P�U`�?Ϳ�r�>Z�
��	�?�7L���.?l����3�?h�6�7?����U?
uD����?O�&�zH�?�Ǿ��?������\_��(�?��=��/P?T�y�v�?�f���U�.<��u>?�f?���?ɻ�=l��>�������?gU�>��?���=V�=�K�>�Ѳ?��C��Ρ�VĈ��ZE?�gJ�m�.�� ��l��@)#�>PO�?N3ھd-Ƚ���>���?$잿�|��.�?3��?����^�(��#�DY�?N��@h����?෡>g�&����?=�,?�QU@Ւ"@m/@sg/?
@�?�?	kɼ��<���^>K8/?�`���:� ���v?�gi?ȏ��w>���0?��A�%��?�`�U�?l�?��j=�yw=d)��F����.`=C*�>��E?!fk��������B��?g,E��&����ž�I�?r7��.�پK7�p��>�������ل��k�>��v���Ⱦ)v9���A��"+���پ��x)?��-��J�r=d뾎=���b�D��>����b���w?�<k����7�3��+�?gG ��B\@�M���?�x���s���"����=��Ǿ�놾?�	�G)W>t%�g�"����0��m�^�f�o�g�h�:��)?���<���n�`���{��:?�j����6=�JU�L�>��c�y�@������?���="�@Ш��'M�?���i�?q��Z�,>{��y�����>yξ�Kľ���yp?Sg?%��>Z=?�e?rü?ӽ��"@!^Y��1?�U�fS��ȍ?u�Ǿa�6>�l
�X	ܾ|����6�>��/��O�w�M�x�)�2�.�>�ʢ=����>���)���_����ZG��;ᾁ��?�A�����̍?<.0��:�����{-z?ٙ^�JMZ��|<8��?�8��i�]>�P���z?�>վns?� ��B�>�Ⱦ��?���;3�?���?��L@͕@��?Ql�@>�h@��@JA�>�1;@�U��5�ȕ@[�i?q�:?���}��%ڞ�t�a�I���[w��J`�I`��� ��'?䱫>�v?��r��?�f�?�t]?�R�֙ݾΞ?p�>N������ƾj�@RG����?e���?X��{T�?l*@�"�?��??T�?��?�w�?Y�k?���	�
H`=r�Ľ�:?tῌ��>��U�%�?�����>�K?~��#������v?i�*�����y�9�}7� ���3 ���	>B;�=uMk��C��%�(�/f&� �｛gھ�A�>GIa���)>�'w�gu�>!����?p�����e>.� ���?�j3���=�!d��v?az��]w�'�r��ۇ>)>����I��oV�O_R�+zG����Co辛�J��0�>�S���<�,���S�����о<f-��������=�9��>S��o
�1�>�Eվ1��?�{̾��F?�K�?�@E�N�F��>�C#�f��S��e�ξ��}��!��$?�A�?�V�Z�i?��k��~�?��?��?�H�>��5?:x�?�K >�W_��Nm�~�V?���<�ℿ��� {��B�=����a?[>+�2}?ߚ��z�?�H��յǽ�y�|k/��-���=>h��@S�c鞿��"���f������i��љ?���?��?`��>L�9@��>I�K�����G6���_�����ʆ�����̾����S�?@�?�f>��A����Մ�7e>��.����>8Fm��٦�;;��@%���﬿��^� ��?*����-���y7���)?��>#���6�]�Ͻ�3����wh�:��3�N��]?�Z9�BUʿ^��uW�>4�W�������8�\�?��e���Ǿ��G�g�3@_�?�Tܾ�(0��
?O��=K�u�x������?�?��++?ǴO��P:?��P�/��?㓐?��=���>�>�>��X?ƁF��a����N��%>�8���?G�_�?�F��|�,=��b�\�?K��� վ�A��Ӑ�6q���@��uʾ���kr<�����=�C�w"@?/1辣��= '	�q>9?�r�� $�]Wz>��>S!��4�f��I�Q�=Y
˾��v?�;@=?����?�<ݛ#@2@��?L<b��(�?�8�΋ @�t@���>�^��WN��Ϙ�<?�վ�j>�s����?m��?�I���DH@����q�@��?Ƕż�1���@�G^>���>Qx�r�>�����=��(���o?
����T۾����<KCf��`���D�����>	 �>Kĉ��]���H�>�����~���ɽ�`;�=�?�>ሉ>��H?��=r�ɽk��j�>@U^?U���?;U�=�]?>��S�}?�?���=7��a>��-��&�K�>35���;����l$�?\W��yWF=�V�:G�>��x�c �dFX<�ƾr������=c�B<6���i�>D�y�O>r㖿�K�>�白lwK?��$>��>��>7P>�;\?9�?6Mz>G~v>(�Q?�?��`>�O�>*��?#}=?�
?�"���߾DϾ�w��(@�?�Q�>�ϯ? ~��誧?e��<d�?��?t�H=�z�{��M=?�1W?��?�%��G��?I�'�Ľ4�I~�����>Aa��Q����{ <��Q��.���'�w�o�~���Su(��]�An��~Ա��ߜ�N�� 0�Qx��E�8>�z>������!�o2��-R������#�b��>�p�����ǅc�sa�>������v?�/7�S߇���{��"P�^;�?-h޾��?��>�?w�B�&��?��?U��?;1D���������Ӟ�?�b���ob�[�R�b6�?� B��Ը��*'?�����b�g��dy>/�v��%|�@c�������*��7��b�C����GJw�=�ƿ����T��#�c���o�����=�p����9�V�1엿��.���=��\�~ɶ�o.�Ŝ?u�S����!��?3�
?��?pr�?&~"���t?&���)?�Y���?�x���w��q��>��@�㏾�a����޿�*��.���8?��>�p�?W�@W��?B5m?a�2?�@�P?��{���=HZM@#պ?�?L��?�a3@ֹ@j��K�=��	��K�8�Z���e?�!)>6���q�@me澊��>�X�>�� @{�?�Te�KM�>'
�?{��$��(��
?������j��>Q;y���?�.$�/*�?����t�?4�H�>�=?�	>�C�>s��<�F�=��=	�?#�z��F���Lm��۲?�x��ɂ��W��V�?��.��U��'�T7?��l����˾���D�����/�־�y�����r�Ts��{M��q�˾�й>N����1���
���"?3�g�]���(j�0�>Nq���PR���
��nu?O�	�ꢄ����?$G����{?o���q�C?����zP���� ��>'ˢ�I�?�]�?�/�<H!t>lʾ���?��
@�愿�\b�����+կ�X���H��+��������<�o�?��@����>mg�����>���L����x�>����.�=�$�rae? ����tB�?C6��{�?QsM�S�%?��Q���?�Ap����?�6��)�?��P�ZH0?>~u����>����U���>@��>0ԅ?^�V?���@��?갘��l�>��˿���?�h��|w���UD@���?}�?P����ۇ�h�NY�?D+�?�S?eL�	�Z?}��H�;+"�ʂ�?	�ھ����y�Ǿ�Oz>v��`����>��<�x�j�#v3���=v�~T����>�!?�?{��� ��̱??�j�(�2�������?���m�?cRj�)@p�?(;3?+��=�� �8��׃�?�*�?<�¼E����>OvR�٤?��v���8?���L �.Ac?j�?���(@";�?W�����?��?3�����>����v���w-�P�������F��=?�(����C��L?�3�?$��>&Z����>��?-��<d���k�龫/?�1�}��&�Y����?w�9?a!?~��:s#T?Ex�3�������>�=ף���,��|���>e�W>�>���HE?�ϕ�E���v�<��fȾ��t����SX�&�9��8�3�=�v?��G���>�!?F�&���<�N�6���K�W���?N�F�i|
?�7��^3?��I�riN>�6�"�=����M'r�����F���/'�?,�ʭN�N��'P�����Zy�?��?<�>Z��>�����x��v�F�C�뇿�$���'���3=��^��bb>M�@��䱿��n>�V�,ؾWW���D0?����bb�=��>��?��ͽ�.�?���?��&?zㇿbH�Q�?�2�?ng~�e��g��>�#C�`�<�o����1�[�o��>�[��	I���ھ���=�ž���;s>��=�����k���侢��>�_K�z�[��U\����>�E�������C>?�ؾ$��>J���1�<��ƾ��5��6=}))�Q�G����7�+>�+��	���'C�M�>��0>)�V?���>��-?�0�>��������(y����U��>o
p�)�_�`�.�;d��Dܽ�U?%�S=��+>tr>D&�?��?叾O?J췼Ai�?@"�>0�i>O(X�%��>C��>򓀾/����H$��D�?
Y�r��>�V.�α�?�{K>Օ$?����.?���>\����̤>@�˾)�u?3y��&��=�P�>��y?sS�>� ~���>�B����)X�>�p`?o|�>w�>�K�>�k�?��?P�?d�������@?3@5?��b>�S�<M%P? /?����Ql���:�u\�Qa���ֿso���\����a��PR+�(AS��$b�f)�s,���K:?PI�a#���$�r��=����~���9�΅=Z@�f�H?5;P��EC>���=�?�)_>U���N�<hs#>�D'�w6�;��T?c�&�c�*?�\������b�k�(�	�Uю� ���?H����������龧b�>iK��A?���=թ���Ǆ?Ȁ	������? #j��A*?��>TRL�b#���+>l�k?U�ܾ2i�<ڨ>i/?���>�iQ?�$>���>o��>�F?=�=�J1;��L��*?��&�w�="ֿ�k�?u�=s�k>s:D?��?��T?ߧ�>����u�T?	�>�U��=��8�V?)G��y��ax?Y�<��"�?>�^�"�?nPX��1>�>Mԗ=�5��U��gŁ���5��&_a��Á���?�?%�+�J�+�����>:3/�	�1?R˧=1�z>nTf�sl���1ӯ��ܠ��A��s���'󄽠l[?�������u��@��>���`5��>�پ��\?-�?�ľ��1?�g@�Y�?[R�>�]?I� @pE?��H?�H? L?���?�c?�4�S�?}�]�A���P�6#;>$Y��X�Ɇ�>]�w?��s��Z�@ӟH>oL�?
Q3�L��?,�!�l�I>�<_?�G�?��
���Z?h�?I�e@}��?z�@�q�<�DH?�ز����=���lx>�	?�K@w ���"@1w��� ?G4ȿ{y$��vx>�E�>뤍?��O?�T��zN=#D��=�S�AN@�����?hrF?ꢄ����>�ך?��@���?���?'\�?��@�f@�� @`3@c��������8?S4@%/>ם7>�v�>��@`���Q�? :@̎?���U4U�e�@�Z?�"�ΰ<��	s?�@3>S~�<ߩ��5t?���~�->���;3=xo�>�rW>̪S��H� !|?��k����>3>���L?���>�r����xc_���?;+�?R�*?�
�>(�@��v?��H?7?�>��?~��>y�E?�Y >���?�"?��>���>0�?�Z�&V�l0���8�>JPJ��F�=/�p�s�lCþ��x?s9c?F<��,��9����E?����O+�>��?7��>N�	��̒>��T=�ܒ�pݦ=ݼ���>? ��>�T?��Ծ}L2>s��=���=����$�j\��?9��+�LMB��>ʽP�=K�]>{�O�]묾{�=YJ���
?�Ҋ��)�>*� ���KԾ��@]���>�@�$x���g@����(3����9>�Ӎ���"�������F����?R�?�O�@�:b?�69����ʞ�!�U?6�ܽ��W��WK��w�>��վ	�>� �]�J����U�5�O���<��Z=�ñM���8��f���G��OO���M��υ���ﾒ
�V$?`����=�Vn?��;?L�M�ЙC����>'��>�>��H?�ԝ����QM��&_��=@���O���숿
ɖ��征ۣ�m��?J��?�>�@��q��
}C?/o�?����[�?�	��;����퉿|>$ҙ��U��[��7�>����������Ě�>ӎ��	XO?����"��.;���o�?sOl�`�Ͼ��l��Ľ?L"=�v�:X���?~����7t������?�������Z�=�$?�炿	�����Q��Λ�j��\�>≯���>�z>r��v��O�T>��=W�4�"�v?t\x?`r����m��`6?���>�8,?)EI�)��>4�ƽ��?�p���z����ᾄc���B+����=�=�Ly>�e��a!?�d�����N1?��q3��k5?�������r�>���<�h�=�3��2������&��N���z	�}๾��>�MϾ�<=*�{��{�>eO�4Qc��U������?\L;�M4D?��A��7ɾ�rf�5b�?�K��Zf>Hn�������8Y�R$��J1?q�>���[y'?�	�@HD@�_����U�S{�>�>l=�8�>N�?�w`��\�?0�?h?������5>�?�ֶ>�
���D�>ה=?��y> ,�*!>���?y1�>l���eY�=OO?�fN?c>ҿ�b�?,q0?]/���2��3�K^?:M�A%�Ҏ��U���>�  �	]���
��v�H?��M?�8l?�|=?�Dh?	@z?6%%>Ń=>̉%�)��"��>�⬿�����>�1ξgо��B?iS��9_��S ���L?C��<�7�X�G�M�U��N���a�>�1��>�+��"�>��"�K8�=�<����+?'�3>=�¿�R-��?��&�o�+��>�ҵ>�靾y�<����?�?GD���ʾ�a;?�[�?����U��?�����)�?p#���E��ܽ�H��ٌ����1�����LD��B��P{�n,?�"���?�gL?�a#�6�A?°ݾ�,?����E�>������>�D���_?��)�R�a?N����;R����?�0��-?������L �0�\�������ᦔ��J�d�پ؅�����=Pgn�����q(��A�7>����K{���u(��3��>��
?�J�?����h�/@ٱ�?wz�1a��ߑ���־
���s�1��g'�91�d���@��� 3@�_?NW�>�@���F ?�����������
��?�G� x>ɡU�lt�?������)���Iw�>%ǿUb��o�R����r���&���i�pO���ê���g��2����?����a��x���$}�Y����D ��ٙ��@���⚿�߾oxĿb��9�?H����L"?�?�-����v?�Ɓ���y@&����;�?@؞�`W��	,
?:?ϸ>�ܳ?>�0���#@'�a?C�?!�?$�9�:X>�e��;�o�?y�>�P�� �����?��uv�>�^.��x�>>N,������f����> �ž�� ����>��.�]ǡ>�9E����>_
��`��>�·���k>\8e���?��þ)#?o�����?����sS�>J�&��]��?|d���Ƹ>�0S�?5	�'��>n��7�*?�.?��=K��43��*_�?@�?�o��{��<UTa���b?eEI�!w>�^_�و�>� )�l�߾�in�n.�>;־�#�vxt�Y�n�f��_O��mJ��7���a�=���]�g{����c��8D�1`����Q�/�ZY��!�aľxM�Q��>����[>��"�bf�>��Ӿ�\4@*Y����>v^ӿ� ���>]=�y����0b��ه>&�j�d�?h��?X!�=Ѕ���<�=V����P_��7�N�=;_
�F K�c�����/?��۾޸�˝?v?ĖѾSW�j�-�o��? �������;�_?�`ž= ٿ��~���W�'���r�|w>��Կ�L=.C�F����`��Z��>��?����	ſ��->�>#���:*��&�?]�G@���>"G?��_:-�U@��w�
u?��߿��?�Ȫ�("?OF�>��>��{��l?i�,��,?��ο���@}'�=��@�$�U�3@՟ �I�0@?��>�H	@23?��@ �f��|>���S�@�?��t9-?�|��3�@�Ǿ�?`�J���?b�j�@Û��h���`�?d�8���H>h���n�@f�� �G?HٿBd
@���Q@}�#�X��@]�G@���0{���C=��t�ݻ?P�a���?Cھ5?���d`��>�J�=�A��)�F�?T�
?�e�޾ôV����?E�>�=�$�k��?ϵY��7ѿ��F���?�'��`�c�LR�>uA@��lj��V�,8Y��A*�v.W�K�)��K������>�{+�<�W��Ua?�؈�Ĝ6�uT|�<Yp? 
n����� ^c��1?��j���v?fC�?(���l�[?1!A�	�@j	N��:�??틿���?��o�hʳ?�ر?����<�=� � �m?X��?YE��� ������?ceh�'�I?`�Dė;������Ѽ����?I/쾀n��II<�_5?(W-��-E������>���"[e��Y�쓿�^�n�5��rW��z�{P8�Q�:��pBi��塽CX<�`>�s��_�Q��
>� U�������~�i������$R-=$~����>�����AQ>���������9�/>ly��QU�{����~Ӓ�gʚ=km��ps�>�5��^|??-_��ߥ>q[����w>���e�G��]���$>�wB��t*�P�|�V*���[�7��>�M����?y?l�>�	?c�p��G?��t�B�k��'���{x>�x��4��T�T�@?�l�ec�������t?�j��1��?��<`a(���?�۝�du�>\-���c0�w$����"�ө���s�?���? ���k}y>(��>?֣?�J@^և�/�����u"ʿ�����>�Y-�T����ⷿ4�������ȟ>�b������r�G��?S>��پY]��]��?Z|�@���k<n�x]����2n?����
�?_1���x�?#����?C��h4�?�����>�h�dv�<�����U��6�Y��?´A��y���I���ߊL�ʓL>��!��cƾ:�������c=9�j���	�?���[,P��y�>#�>�Z��u�g���>�e.>b�?E���p�<T,>���?x������?��ž��?i��[�!@��?7�g@�9 @�#@v�@?"`@�O�??��?P��?'��?�n:>Hi�7�޿�Ǿ�5��O=H)�5��.��?.�?S5�Y$@��>�>5�~
�=�v��_�[�ا>�?�|���=
>ߠžb�p�>0=�>��Q�G��N=8?�!#?o�?�O >g��RZ�}��D���VH�!�>�L��>����Y�?O�0����;�辫W'��:��4���^��#(�>8���"�;�8"�[��>[�>_�=�E-���>�7��G�>t-�?�q�>}s#>�g1>�X�=��'=ڌ�>2!ʽ�� ��D�?��(�}#��c��?z�v�6|t?��C=�Q�?*q!����?��F��E�9�F�]��e��=�d)?r��?�w?�>�>M;�?�>&ݰ�Y�?�ҹ?�?�ȵ����� Y?=o��n�Y�����>��辝r-�Ǩ��������@�y>3��g׾��6�[ň��k�������q�ڔ�VƾL?��:��JP��Q��8]5�,c�E�	>m����k�<|��ﶥ�TWZ>��?�����>1�^�b�?0�o��[�>��F���>>��V>s�>xA��n����`?���?�t�#���J7d����>�����ؾ�����_�>֩��Y��[���7� ��o��M��D�.�1��}MS��ɪ�|�E�����`C���N�I��8�A�)��6�M)�%3?́1�w��?��龋ރ?�`��j!�?����,I6?����?Ԧͽ���>Қ��+]W���u���>-@^?��/�f? �7��<?�Y�U�E?@MI?��>��,��}�7��>>����QOM��W=<4�b��.ž��$�ꨀ���>���l'��Fܾ�/����I櫾Ss��Yo�����>�;�=>��j�aq'?��3�m����mϿ�4�O�N��̾޽h��?)u�=�s�>��g> z?Df�>�Kz>�G�� �u?��<��� ��>k��?`��>�/t@o�X?Kt@��??�>Ɩ�?W@����:��hھ�(�?͞�Y꠿���+%>"Tѿ��?jI�?��>8Un�'�\>���?�?�Z�>&�??taR>6b�?+
?��?G^?d�@���?��?O�?�?5̷>�ھńY?v��>[Pa?�������?���?�y3?��>�f�? �4?�>�>�����>[x?�p��U��6��1'?�1� �T���9��c;�L��y�d�d��P�=��u�?��?_����ӿ��E�:C��(�տ��ʾ>��=a?�
���v=�A�?y��?8��u�e>'��?5V?!��Ԯ>�[?4ԗ>���o+>*����
��&�6i�>��}=���������<�m��X��D�?vȿ���~(2?�f ?�п$�0?ޝ�?�Q@�'��o,@���>�j�?+�8�<ጾ�<� A?���� �?jCξ��?�%���3��x���+�̟���� ��և�Z�8�s��m���"���?Q_�^=#���5?�+�>��]>�LȾ�%�>\v?�S?�;2����#
?[�?	y �*�$>��?/��?^�.�hﾾ�)R�E���N�?�	臿?�Z���>◐�nQ>N����>?���� ���^]����� ؾꢄ�?�l�z`?�h�?L���(>1dF�|u?t೾�/(?)��L>���ɐ��T�2 @��ÿ������7?��@��Ͼ],���?s�ξ%e���cI���º3�HՋ��C���>�n�?z��>' �?�,d?�i%@y*?�H@�&�;���?�džъ?��[�Ͻ?�@��Ƃ?�r
�!��>�4�=d@��?EU?�Ak>��?UH����H�*��ꢄ�{B�	6@����x3@����B��?"�o���[>�þY�-?YR�m+<��4�?`�5>o���-�4�	���U?Lb����?y�,�c�?�r�?�V�?�@�����?��?@�?��H���a?7��?��?�ZM���?������X?y���.@@jǹ���*@Q%���@9������?���?�S��+ϋ�P�?��?���?���UZ�>�(�?K��?F����8E>h;ľ7Y���@	}8��?�?w3?RD�@o�<
��?�@�>�_�@�?�A�?>���ْ=���<�.����!��T�?�n���N&@��\?��?�×?:�@�n>�?ْ<���?)&y��<f@R�B=fT3��
��ի?{�c?+aE?&3?��?�s#@��d@��@8��?�'@Q�@��??�3b?1c���?@*jx�Ok/@���crq?�A�?�R/@�c�>��?��>�ɽ�/>�+���d�L�E?8�����x��<*Z>����@-S@���>ܟ`����>�ֽ>��?��?^�K�����X���T?m��>���?@eʿ���? y�>�@?����2>;B⾏��>��ο�q(?ǜ��;�z?p�ſ���>06���DD>�m龲�1>���J	G?9ݤ�&���ӫ���h�?9�e>���=8�;�s��?�vu?��.>��]�w �>���>���_�<�j���
��͕?0>0�P�?#!�6}I?��=�ۨ�?�R�?�->��g��M\���?��?0>^Z;�䗿�[4����<?+�>��a��n��R��򬫾��-�JxZ>��F?�B�SM?B�\�4��>�ǿ﬒�������|<�`��$P>:��P�9?�S���?ᘋ�>�'>\��?��>R�p>��K�.U?)m�=	�����t�1.�c�f:�B\@#��ڦ>'>Җ�<o[|?�<=ʃ?�a>q'k?(>�:?,?>ן=�鋽u��W��>��m?� �+�R�R,�N�>ϩ����돾�? �px?���iþ�k)?=�P���
Z=�ms���s>� ��p�w=��j?��=`�>��2>��s�A�>��}>1�=S.ɾ��f?��>*sV?[D���>�� ?��
?��վ�c6���?[겾�
?f��ؼ�T��sӺ�W�>Bs?U�!?�W>�
�>�!�>(�?F��?P�+���q����;�!�V�;�u	��8� �F��>��4?I�%��~~�T�ݾ�� ?8(ԽC�����X� ?� ^��3o�J��J"�>4��yj�a����v��,���죽����T��y����Ͻ���ـ�1���f=��ݾ�؃�Ȭ����$?�_��W`��W_>�:?��$=w6�;���>��˾��߾�+�>	����h�>/���C�?�V��F�d?3�?��>�d�>z#�"��=�r�>i;{�4AC@M!�?%��?�>>��E��y=��>��1|�`�¿��?�f��{�.�B�ӿ�j̾kB�=k�ž,�c��?�w;?��<�s��D�>��^?�ｾN ���`���<��gv����"��R߼��>��?r���S�?%��KF[?�� ��.�?!����l�?��(>�;?<��6"��u����>ZJ���I���:���A}?�
 ?Hb�?\%O?YF���&���>��꾷��Y��?�����OD����M��?*�d?���<��=@�/�?g�c?���I��?� ?g�>"0^�E�>��M>N%>�i/>X�����[�"�e�=v�o>t����O�!]d?7�� S���1Y�c�i?��<ٿÿ�r���v?O����?o\�����>(Ѹ?�9�}�?1W??�0�?T�>�s�?~�?��y=����1ξ�l-��q���L���� 4����>[h�?A#��)\Ѿ:_�=@O�>K����m`��J�=uŅ>�N��$��>=��=�2��L�c8����^>�$?�L�=X��> oH>��
?��?�o�?�.���?̀����?mM���?t%v?��?����O��~���R��sS�>���?��ܿ�\0?��M�ٶ�<rw���������*��I��e%�>���>f�ؾB!�LHC��6A?��?%ދ����<ࢿJ߼��`?���?[�W�w����^�yɋ�b����1*z�)�A���i����>� L�mʠ>:�Q��?��:��нZ�6�hڷ=�n���+�>&�ϛ־ӹ�s��[,���=�"F�sU)�^�g���ݾ�D����ջ\���H?~Y@�<ѿ�]�>5��ǫ�>�!����������_>M�Ҿ���>(z�>"qi��=�m���-�<vY�>�A��g)����+����ԓǾf]�?0��>�)}��(�t~?�?�?/�����{�]��?m�B�K����0�#�S?/����m='��� $>�쀿�v��v���ο�LZ�֏�?+�z�J�ʿ�cv��ɷ?K ����տ%���	�@&⍿�~'��3c��
?�oS?_��:nȽ�������Ä��ײ���0u7��@͝�`;����z��羾��x��4t�|�w?E�&�fM?�^���\�L(���� �����Q�[�9�ǿ'�Ŀ�I��k`����ҿm��e�z����=sҮ�_c�=�/a��ξ�}�4�">E3I�'u?U0)����?�$�E�<�a��\�?��Z����>)x�����?y����t?~8���X@��U���H?�c�?ګ����>*ZJ�Ӄ�>�?Ň�>-X�,>	��[�`�R�`��.�>ִp>_ǽ�$���GX?� �����m�?������a��������0P��`�i8���þa�����T�w�+=�IZ?t
�?[��>),���������?�h����z��"��x#���V���v�@����?�K���@mv��C�=�L��h@	@�nr=w6�;��s?
T��篾��/��h���v~?[*�ߤ�?I���\��?��5�����zf��IU������"��c,@� �?Z%>>0�?�,��Т���J�}�ƾ%�h��Ϣ�v��y@�����?1�����&@ٲ�[��?�&�ɚ�>gZ=���|3L�3f��/W�r{�4Zt�wM	>�O�L�I?X�����%>�Y�>B?�k���י�y��9��><����
?e��?��O�J�B=�������0Ѿ�ꙿ��&?���v"=-��뿒���{�=��>39G���ſ�!>���?� �Fxھ�f
?���?@=?^��?��_@��w�?)@D��?M%�"��<��?�*x?�Ჾ!�r?%�>�g�>�M���=�I�פ����x���>-����`�UNF����>�`6���:���;�L�	�e���C�����饿�6��ꢄ���?�l��L��>�W���?�L�¾�.?��Q���u>�Z�3��;���s��8�>2��=�'��+)�>�4'�c��>��%�^m?�;�ѫ�pG@�a�n>옿�$��1Jپ�+?�d�;�,�?+0���r�?� ���?�l��R��=�(1��?�X��_־C�n���?� �M�� 2y�s�?����#��71m�?
?F���oU��z� �G?�$v���v?ӨԽ���>�>H�o�9s�bF���_��G�\E�g�o�Ї���%>��e>��u���G�=I���>��>ڙ�jd�=$�K���?�Wp�-D?��y=3G=�]>�?gc&��|<�҇˾ke??�0H�Nɢ��_X�@�?����^>��
�n?ݙ;2B���6��}��$��Z����[H?���d]x��-|>�`����}�Ӿ�N�>��D�w6�;3��-�f��Bȼ)x����n�:'v��Ե�}@��#��X�>pB��;����8�����=+�W��$���U���@��G?i�.?�s?� =�f���?P��e�l��?�ܖ���t�Lߐ�CQʿU��I��;B߆�RR�<Ž�>�?i����?4�?���?�C>B��?��g�&3@�Ӿ�$@�e<�6?�)�p�r>����]���;��Zؿ>?��ꢄ��]?}�۾��ݿ*�p�A����v>Vɛ=Ɔ ����|>��B��A�Q�g�"?����u?Xf��1��K��=7?5^R��B�?�3��'�rk<>��|�I�N�.�ѿ������=�撿�B?�x#�8�@�+��d�>~��!�<÷S��V?������? ���9�=��4�JB���J0����?�]�[+?O�ƾV�>|�*�DQ���2�r�?�/��4`��"�j�1?�b������5�>�@*�#�>��K���>S���)?�??�N-�7p����=� N��>�Mr���+���?��=��?Ή������~"���@&7��F�?������?���{�>�"$���
�WȾQ���+����Y���>̰ﾲ�;&0ž���>�{-?��w��
=x{ھ�'?�E�C?w���� �=I࿄9�>��g�������>� Q��A@�B=?-J@{�¾8����|���gξd���j��Z�������M�?���?�՗�w��G����m?�$f��f<x�8�MJ6��c����<���5>Y�s?Ԟ׾ָ
@\I�?jn@�FB?K&J@�?Ϫ�?����),�?�Y����p��������>k�;>ј0>�=�?�2�?h~> f�?@��>;��=h;I�˺=
i?;?[Ҿt̼��,?+=�?w6�;<M�?���uCc�*O�mп�)�/O
��BY��M�z�����,���*�R���~ >?X��������7�$�\?��C��	Z�V�묫?��#�4��?8�|���|@�1����;@%QX�ř�?�x)�<L�>�� �?��e�d��?�y�o���u����(��k��wN�*a��])@�)��Џ���~~�eU@qE>�T���UA����?�6�ǆ��p=��
?��?�����[������ƽ� ����Z�*����'H�J�[��կ?� �?ｔ?�#g�B�4���7�틛��V;��m�?���A���س�xJ�?d{�>n�f�_�k�c��?ؙ8��'���lu�>ȝc�;��?���@<�_ك?e[Ҿ���?�'�ɒ�?|�1�>��@z:�7?�?x�l���R`��Q@��'��_�o�U>$@f�g�tZ��M�h;ľM����p�?���?x�1?
$�Q��>G�-=��ž׽�����:�Y�A,D���?�@�:'��%Q>��.?�����Q �>��s>��=�I��VF?������D?��F�aL�?�(�?M4@X��?��L@��@O7@sW�����?��I�J�>{V����V>cG2?���?|v?�/�>�}6?���'%����>��C����8�=6���`
?>����YD?,^�<�
?DE?��%��ሼ�����[�>�#���!�>!}��wn>���>IP?�3�=a@羘^�>�
��X�?��t�4��!���5+?�d뾼�>����YU)>&�=? ?�\���Ű>�þB/�>9���/�?0��Y��=A5���2�?�B+�Y;�>S��ֹ�?�=��T��q�G������{�C4@��n����о��C�/���S���ϖ����[���
?:��>�s0�. ���=��z;?ߍD���w?h�Y���g?��C��=�{d=�}%?�&+�N>̾�ƒ��	>��/�����q�q�o?��P�v^�>K	��F�?� *���>��5�yj���X�\�=�QB�� ��6�J���>�����=Rw\�U�V?�T1�������@x?�r��c&�MzY�2a??�&j��Ϗ�2�辂��>\X��"a���E�ȥ5?S�x��\4@��;��_�>�����a�GԦ�U�	�[$��H�1:�&�0J��M�?ɱ�?��9��v����=�1���ۆ��覾6AZ?�R�a���>t�#@��ƽ�.��	N=oR�?f7=\a��2�n?���?�ާ��z�b��?::>{������J�_�@���.��˽>p���R�A��_M?�?>��'%Ⱦ٪/@`��>f�q?/�1@,��?^�ֿ�y�?��v?���>7�׾,û��@6��R}��a�>������RԾІ&�C�8?�<?�����D��ˊ*?Û�>2k�>�c�ڂ>��]�N���ľ:!z?�XN?�'U<$�d?�։=v�p_���}Ľ��4�[��_��Z�3�Ou����E#�B�=�6��1�>$b��\T?�,��@A�ş������y󾥂�g4�1Y��4����m,��/Ǿ��پX�>��2��
?�Wc>b�I�Q웾�0о*��?�����?�\���?h����SO�ϱ༜��>m�w�Ş�>U�(��� ?wAP��Ph���@]p?P�N����������?pC�!�{�ߝj�Q@�>�w��0�>�J�<�8�	�7�q��=�-Z��h����_��4y��7Y��#��}W���>��#�BMj�86]���>~\�R
a�L����@?� ��NW*�Vߪ�m�&?v���sS�>���%�>��g?�s�bb�0ΐ�^�>d��끮��Wr�#��XZ �[<���� ?��E>E�?�WE?g�?�GI?���3G�>d��=w�3��:���>Ȗ�8�K�����U5��,˃�ɭ��I��̿|����9�I��ݦ�6����t7?�y����*>@+���?��>�}y>x�f���?e�>�><b����?�&�?ň���<��?\��ꢄ���?�ؿ;����w��dw>�v��⃿�jU������6m�#(�?�T�?�v)>��Z�h��>/(ü�k�?{b�ׇ�*�e����
�π�>��L�Z�������aI?�i��J��4]ܾz�N?ZQ:��g?`��8*�C-��U��)��X?ǀ�>X�K>�w�Р?͔}�m�>���%Ǿj��>>ϹJ��Be>h*���R?��v��! ��K�1��?��?��/�2]@��@Qώ��ʼ?�fN�XX,��d��ؗ>��v�F�w�!�����+@Q\� ��@�3�?{�*���w?y�@���>��߼п>�����?X;�>/�ZU�~f?�K�������?��>:��F���R�U<C��-?1���������nǾ_��>	���b���=����'�z�,��*]7>��+��{3��+�� _��}g�p�y���r��Λ�-e�0�N?���>/X>5�%=R�>,����T�L�ǽB5C�/�?)s?�o8>ڟw>ֿ�=�2�>V�P?m�� ��:?�>'�H>�QU�ʖ>����󾗖Q�|>
?M�޾��'�J
̾j��G��y�S>Vaľz�+�Q�Y���^�ķ�)����>V�˾��
> _'?�@?��?1�`?�?��@?2�E?�H�>IԐ��].� h����8�sS�>����9%�?���[���ti�l�����x������l�4K�����z���=�U轛o��8�_�n��L\u� ��I��'��cM�2}�?�n�vڨ?�%Q��C@.�־*N@�n�>�[-@e���J<4'���?��&+�X1�����>u�����+�IV�?T��>�@��Ze�?4Ƚ� ��A�A�l���H�����K����?Ȳ��I��$!P��
?�E>,<ѽT����ŝ���j=�����*?�a�� �>j�}�:Lp���p���������G�>QM����wv|���r>�a���:�?/�u�A�?��n��a>��-�	�^�6�o�]�B��S����R���G��ž�
x�	[G�MM_�m���fn�����(9d�Fd��ɘ����?�w��t:�-�9�|,e?��g�7���CI�'S�?�R�}ɧ�]�;�%B�?�ɾsS�>V��?J�ɿ��?�G����?֯�Ԝ{�k m�"�>GX�/ŕ?�z�?�$��r&���C�>uq�?���?]Yy��O<<RB��F�=�08�=&@릠�����	� ��ȗ?ղ|��ݿ;����M�?"��n�?�ن�ÿe?L79��7��.UD����B@��%��0�X�����w��b��
ϟ�N�տ�<���b���_���?����o�>5���< ߾Pf��� �1�(�`�B?p�>ӻ?A�@-�?:�H?���-��?RI��hG@��@̉?L�?���["9���>���wm����_?0�=�������}�¾Lbſ����c�?h�����O�0�^<��1@Ƭ�?!)?�@Nů?���>s׿օ&�2��=�>;x��=��=�}+>�	E>S8�=GuT?Xŷ>�I@�)?+Ce@�N;>S�?e��?S�-;}� �O8�����>��i�p����H?��Cz�0���&R��kJ����P��Em�������xT�5_?je߾|о=І���;��Mu��\�?3|�V�տ�IP=7)�?�D�}���M�;���?�p��%w����>��?$M��ǒ��TM��ч>U�D�X��=Z����
�>M8��O�?�c�^�R����Σ�??����.����>!�>)ܾ6���!־�|�?Z��>B�ɿUq�=b���U?s�d�a�=���#��?�h�}�?��¾ͧ?�g����Y>��q>����M�=w˓�o�\���!?Aq��聿8p�8f-?�P�����]��-�c?J�=�����b"�B�?��E�Y�r>���Ɋ?&���G?J"˾�2j?-=پ��?M/����?�Y���}�?y�7��j&?��|<�Ƒ?G��{(w����=�#g�*h���c��Y�9.?��C��U��F,���?�H��^�(�!?��+�y&S?��|���9?,���]p�?�6�?����w����ﾕ"�ܐ�>���ꌾ�NɾFF~?�{P��{E��1�v�l�F��Xx�8 �ӟ>H`~�(Fx��o?�N�*?����B��:վ`�}���\��O�'�=�ՙ�#?l h?j�>F�D�3ث=�?�>}�E��ɘ�6L��Ċf���[������1>[�c��7����?np�?6}3�カ�+�G�k
�)QȾ&:��{���y �����i��5��ߡ�>���=q$½ƛ����
���F����?td��Ų�����@I/�vI�<c����@�`9?i"C?��K@aL����p?8r����?\�ھ{�H?�(V�x|�'��|T?���9�M���r�x�?�KS�gп�V���)�?�Te�J.����Ӽ?@��A
�K�#���v?�A��I��9�:��:��m?�?��,�J�@��%���
@7y�Oqm?ԕo?#$>>{��E!��r��X�?��\����P_����?�5K������O�{h�?��\�u��u�e��!>8�>���8��l>�p8���?S�^���Y=MII��2�?6GB��w�pK���9�?�0����,��G?k�]�f#��ҩ��%8^?:����=��ư�|P�?�� >�?       �t�b�n_samples_fit_�M@�_tree�N�_sklearn_version��1.1.1�ub.